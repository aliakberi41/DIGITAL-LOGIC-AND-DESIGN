<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>56,-4.5</position>
<gparam>LABEL_TEXT D FLIP FLOP</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AE_DFF_LOW</type>
<position>56,-25</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUTINV_0</ID>4 </output>
<output>
<ID>OUT_0</ID>3 </output>
<input>
<ID>clock</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>26.5,-17.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>BB_CLOCK</type>
<position>21.5,-27</position>
<output>
<ID>CLK</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>79,-20.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>80,-28</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-23,40.5,-17.5</points>
<intersection>-23 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-23,53,-23</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-17.5,40.5,-17.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-27,39,-26</points>
<intersection>-27 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-26,53,-26</points>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-27,39,-27</points>
<connection>
<GID>8</GID>
<name>CLK</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-23,68.5,-20.5</points>
<intersection>-23 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-20.5,78,-20.5</points>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-23,68.5,-23</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-28,69,-26</points>
<intersection>-28 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-28,79,-28</points>
<connection>
<GID>12</GID>
<name>N_in0</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>59,-26,69,-26</points>
<connection>
<GID>4</GID>
<name>OUTINV_0</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-6,3.77107e-007,116.4,-60.5</PageViewport>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>54.5,-4</position>
<gparam>LABEL_TEXT JK FLIP FLOP</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>BB_CLOCK</type>
<position>12,-26</position>
<output>
<ID>CLK</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>12.5,-16</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>12.5,-35</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND3</type>
<position>33.5,-17.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>9 </input>
<input>
<ID>IN_2</ID>8 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_AND3</type>
<position>34.5,-34</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>10 </input>
<input>
<ID>IN_2</ID>18 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>34</ID>
<type>AE_OR2</type>
<position>-55,-17.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>BE_NOR2</type>
<position>66.5,-18.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>BE_NOR2</type>
<position>67.5,-34.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>GA_LED</type>
<position>78.5,-18</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>GA_LED</type>
<position>79.5,-35.5</position>
<input>
<ID>N_in0</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-32,23.5,-19.5</points>
<intersection>-32 1</intersection>
<intersection>-26 2</intersection>
<intersection>-19.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23.5,-32,31.5,-32</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-26,23.5,-26</points>
<connection>
<GID>24</GID>
<name>CLK</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>23.5,-19.5,30.5,-19.5</points>
<connection>
<GID>30</GID>
<name>IN_2</name></connection>
<intersection>23.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-17.5,22.5,-16</points>
<intersection>-17.5 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-17.5,30.5,-17.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-16,22.5,-16</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-35,23,-34</points>
<intersection>-35 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-34,31.5,-34</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-35,23,-35</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-42.5,73.5,-30.5</points>
<intersection>-42.5 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-30.5,73.5,-30.5</points>
<intersection>63.5 3</intersection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-42.5,73.5,-42.5</points>
<intersection>31.5 4</intersection>
<intersection>73.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>63.5,-30.5,63.5,-19.5</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>31.5,-42.5,31.5,-36</points>
<connection>
<GID>32</GID>
<name>IN_2</name></connection>
<intersection>-42.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-35.5,74.5,-34.5</points>
<intersection>-35.5 1</intersection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-35.5,78.5,-35.5</points>
<connection>
<GID>42</GID>
<name>N_in0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-34.5,74.5,-34.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-18.5,73.5,-18</points>
<intersection>-18.5 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73.5,-18,77.5,-18</points>
<connection>
<GID>40</GID>
<name>N_in0</name></connection>
<intersection>73.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-18.5,73.5,-18.5</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-35.5,51,-34</points>
<intersection>-35.5 1</intersection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-35.5,64.5,-35.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-34,51,-34</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36.5,-17.5,63.5,-17.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<connection>
<GID>30</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-12,88.5,-12</points>
<intersection>30.5 5</intersection>
<intersection>88.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>88.5,-31.5,88.5,-12</points>
<intersection>-31.5 4</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>64.5,-31.5,88.5,-31.5</points>
<intersection>64.5 6</intersection>
<intersection>88.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>30.5,-15.5,30.5,-12</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-12 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>64.5,-33.5,64.5,-31.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-31.5 4</intersection></vsegment></shape></wire></page 1>
<page 2>
<PageViewport>-9,3.77107e-007,113.4,-60.5</PageViewport>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>54.5,-3.5</position>
<gparam>LABEL_TEXT JOHNSON COUNTER</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>BB_CLOCK</type>
<position>2,-25.5</position>
<output>
<ID>CLK</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_TOGGLE</type>
<position>2,-41.5</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>AE_DFF_LOW</type>
<position>22.5,-26</position>
<input>
<ID>IN_0</ID>33 </input>
<output>
<ID>OUT_0</ID>34 </output>
<input>
<ID>clear</ID>37 </input>
<input>
<ID>clock</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>43</ID>
<type>AE_DFF_LOW</type>
<position>37.5,-26</position>
<input>
<ID>IN_0</ID>34 </input>
<output>
<ID>OUT_0</ID>35 </output>
<input>
<ID>clear</ID>37 </input>
<input>
<ID>clock</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_DFF_LOW</type>
<position>52.5,-25.5</position>
<input>
<ID>IN_0</ID>35 </input>
<output>
<ID>OUT_0</ID>36 </output>
<input>
<ID>clear</ID>37 </input>
<input>
<ID>clock</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>47</ID>
<type>AE_DFF_LOW</type>
<position>67.5,-25</position>
<input>
<ID>IN_0</ID>36 </input>
<output>
<ID>OUTINV_0</ID>33 </output>
<input>
<ID>clear</ID>37 </input>
<input>
<ID>clock</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-36,12.5,-25.5</points>
<intersection>-36 1</intersection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12.5,-36,64.5,-36</points>
<intersection>12.5 0</intersection>
<intersection>19.5 5</intersection>
<intersection>34.5 4</intersection>
<intersection>49.5 7</intersection>
<intersection>64.5 9</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-25.5,12.5,-25.5</points>
<connection>
<GID>19</GID>
<name>CLK</name></connection>
<intersection>12.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>34.5,-36,34.5,-27</points>
<connection>
<GID>43</GID>
<name>clock</name></connection>
<intersection>-36 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>19.5,-36,19.5,-27</points>
<connection>
<GID>39</GID>
<name>clock</name></connection>
<intersection>-36 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>49.5,-36,49.5,-26.5</points>
<connection>
<GID>45</GID>
<name>clock</name></connection>
<intersection>-36 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>64.5,-36,64.5,-26</points>
<connection>
<GID>47</GID>
<name>clock</name></connection>
<intersection>-36 1</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-13.5,70.5,-13.5</points>
<intersection>19.5 4</intersection>
<intersection>70.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>70.5,-26,70.5,-13.5</points>
<connection>
<GID>47</GID>
<name>OUTINV_0</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>19.5,-24,19.5,-13.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>-13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-24,34.5,-24</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-24,45,-23.5</points>
<intersection>-24 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-23.5,49.5,-23.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40.5,-24,45,-24</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-23.5,60,-23</points>
<intersection>-23.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60,-23,64.5,-23</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-23.5,60,-23.5</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-41.5,22.5,-30</points>
<connection>
<GID>39</GID>
<name>clear</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,-41.5,67.5,-41.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>22.5 0</intersection>
<intersection>37.5 6</intersection>
<intersection>52.5 3</intersection>
<intersection>67.5 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>52.5,-41.5,52.5,-29.5</points>
<connection>
<GID>45</GID>
<name>clear</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>67.5,-41.5,67.5,-29</points>
<connection>
<GID>47</GID>
<name>clear</name></connection>
<intersection>-41.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>37.5,-41.5,37.5,-30</points>
<connection>
<GID>43</GID>
<name>clear</name></connection>
<intersection>-41.5 1</intersection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport>
<gate>
<ID>49</ID>
<type>AE_DFF_LOW</type>
<position>27,-25.5</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>40 </output>
<input>
<ID>clear</ID>43 </input>
<input>
<ID>clock</ID>38 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>51</ID>
<type>AE_DFF_LOW</type>
<position>43,-25.5</position>
<input>
<ID>IN_0</ID>40 </input>
<output>
<ID>OUT_0</ID>41 </output>
<input>
<ID>clear</ID>43 </input>
<input>
<ID>clock</ID>38 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>53</ID>
<type>AE_DFF_LOW</type>
<position>57,-25</position>
<input>
<ID>IN_0</ID>41 </input>
<output>
<ID>OUT_0</ID>42 </output>
<input>
<ID>clear</ID>43 </input>
<input>
<ID>clock</ID>38 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>55</ID>
<type>AE_DFF_LOW</type>
<position>73.5,-25</position>
<input>
<ID>IN_0</ID>42 </input>
<output>
<ID>OUT_0</ID>39 </output>
<input>
<ID>clear</ID>43 </input>
<input>
<ID>clock</ID>38 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>54.5,-3.5</position>
<gparam>LABEL_TEXT RING COUNTER</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_TOGGLE</type>
<position>10,-42.5</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>61</ID>
<type>BB_CLOCK</type>
<position>7.5,-31</position>
<output>
<ID>CLK</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>11.5,-34,70.5,-34</points>
<intersection>11.5 6</intersection>
<intersection>24 5</intersection>
<intersection>40 4</intersection>
<intersection>54 8</intersection>
<intersection>70.5 10</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>40,-34,40,-26.5</points>
<connection>
<GID>51</GID>
<name>clock</name></connection>
<intersection>-34 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>24,-34,24,-26.5</points>
<connection>
<GID>49</GID>
<name>clock</name></connection>
<intersection>-34 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>11.5,-34,11.5,-31</points>
<connection>
<GID>61</GID>
<name>CLK</name></connection>
<intersection>-34 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>54,-34,54,-26</points>
<connection>
<GID>53</GID>
<name>clock</name></connection>
<intersection>-34 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>70.5,-34,70.5,-26</points>
<connection>
<GID>55</GID>
<name>clock</name></connection>
<intersection>-34 1</intersection></vsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-16,76.5,-16</points>
<intersection>24 3</intersection>
<intersection>76.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24,-23.5,24,-16</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>-16 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>76.5,-23,76.5,-16</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>-16 1</intersection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-23.5,40,-23.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-23.5,50,-23</points>
<intersection>-23.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-23,54,-23</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-23.5,50,-23.5</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-23,70.5,-23</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-42.5,27,-29.5</points>
<connection>
<GID>49</GID>
<name>clear</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-42.5,73.5,-42.5</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection>
<intersection>43 3</intersection>
<intersection>57 5</intersection>
<intersection>73.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43,-42.5,43,-29.5</points>
<connection>
<GID>51</GID>
<name>clear</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>57,-42.5,57,-29</points>
<connection>
<GID>53</GID>
<name>clear</name></connection>
<intersection>-42.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>73.5,-42.5,73.5,-29</points>
<connection>
<GID>55</GID>
<name>clear</name></connection>
<intersection>-42.5 1</intersection></vsegment></shape></wire></page 3>
<page 4>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>54,-3.5</position>
<gparam>LABEL_TEXT SHIFT RIGHT REGISTER (SISO)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AE_DFF_LOW</type>
<position>27,-23.5</position>
<input>
<ID>IN_0</ID>44 </input>
<output>
<ID>OUT_0</ID>46 </output>
<input>
<ID>clock</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>67</ID>
<type>AE_DFF_LOW</type>
<position>43.5,-22.5</position>
<input>
<ID>IN_0</ID>46 </input>
<output>
<ID>OUT_0</ID>47 </output>
<input>
<ID>clock</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_DFF_LOW</type>
<position>59.5,-23</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>48 </output>
<input>
<ID>clock</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_DFF_LOW</type>
<position>76.5,-23</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>49 </output>
<input>
<ID>clock</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>10,-19.5</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>75</ID>
<type>BB_CLOCK</type>
<position>7.5,-29</position>
<output>
<ID>CLK</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>77</ID>
<type>GA_LED</type>
<position>88.5,-21</position>
<input>
<ID>N_in0</ID>49 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-21.5,18,-19.5</points>
<intersection>-21.5 1</intersection>
<intersection>-19.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-21.5,24,-21.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>18 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-19.5,18,-19.5</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-37,17.5,-29</points>
<intersection>-37 1</intersection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-37,73.5,-37</points>
<intersection>17.5 0</intersection>
<intersection>24 3</intersection>
<intersection>40.5 5</intersection>
<intersection>56.5 7</intersection>
<intersection>73.5 9</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-29,17.5,-29</points>
<connection>
<GID>75</GID>
<name>CLK</name></connection>
<intersection>17.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24,-37,24,-24.5</points>
<connection>
<GID>65</GID>
<name>clock</name></connection>
<intersection>-37 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>40.5,-37,40.5,-23.5</points>
<connection>
<GID>67</GID>
<name>clock</name></connection>
<intersection>-37 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>56.5,-37,56.5,-24</points>
<connection>
<GID>69</GID>
<name>clock</name></connection>
<intersection>-37 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>73.5,-37,73.5,-24</points>
<connection>
<GID>71</GID>
<name>clock</name></connection>
<intersection>-37 1</intersection></vsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-21.5,35,-20.5</points>
<intersection>-21.5 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-20.5,40.5,-20.5</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-21.5,35,-21.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-21,51.5,-20.5</points>
<intersection>-21 1</intersection>
<intersection>-20.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-21,56.5,-21</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-20.5,51.5,-20.5</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>62.5,-21,73.5,-21</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79.5,-21,87.5,-21</points>
<connection>
<GID>77</GID>
<name>N_in0</name></connection>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>0,-6,122.4,-66.5</PageViewport>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>58,-9.5</position>
<gparam>LABEL_TEXT SHIFT LEFT REGISTER (SISO)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_TOGGLE</type>
<position>104,-42.5</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>83</ID>
<type>BB_CLOCK</type>
<position>103,-33</position>
<output>
<ID>CLK</ID>50 </output>
<gparam>angle 180</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>85</ID>
<type>AE_DFF_LOW</type>
<position>84.5,-32.5</position>
<input>
<ID>IN_0</ID>51 </input>
<output>
<ID>OUT_0</ID>52 </output>
<input>
<ID>clock</ID>50 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>87</ID>
<type>AE_DFF_LOW</type>
<position>65,-32</position>
<input>
<ID>IN_0</ID>52 </input>
<output>
<ID>OUT_0</ID>53 </output>
<input>
<ID>clock</ID>50 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>89</ID>
<type>AE_DFF_LOW</type>
<position>45.5,-32</position>
<input>
<ID>IN_0</ID>53 </input>
<output>
<ID>OUT_0</ID>54 </output>
<input>
<ID>clock</ID>50 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_DFF_LOW</type>
<position>25.5,-31.5</position>
<input>
<ID>IN_0</ID>54 </input>
<output>
<ID>OUT_0</ID>55 </output>
<input>
<ID>clock</ID>50 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>93</ID>
<type>GA_LED</type>
<position>9.5,-32</position>
<input>
<ID>N_in1</ID>55 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93,-33,93,-22</points>
<intersection>-33 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-22,93,-22</points>
<intersection>28.5 5</intersection>
<intersection>48.5 6</intersection>
<intersection>68 3</intersection>
<intersection>87.5 7</intersection>
<intersection>93 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93,-33,99,-33</points>
<connection>
<GID>83</GID>
<name>CLK</name></connection>
<intersection>93 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>68,-31,68,-22</points>
<connection>
<GID>87</GID>
<name>clock</name></connection>
<intersection>-22 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>28.5,-30.5,28.5,-22</points>
<connection>
<GID>91</GID>
<name>clock</name></connection>
<intersection>-22 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>48.5,-31,48.5,-22</points>
<connection>
<GID>89</GID>
<name>clock</name></connection>
<intersection>-22 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>87.5,-31.5,87.5,-22</points>
<connection>
<GID>85</GID>
<name>clock</name></connection>
<intersection>-22 1</intersection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>94.5,-42.5,94.5,-34.5</points>
<intersection>-42.5 2</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87.5,-34.5,94.5,-34.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>94.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94.5,-42.5,102,-42.5</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<intersection>94.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-34.5,74.5,-34</points>
<intersection>-34.5 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-34,74.5,-34</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-34.5,81.5,-34.5</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48.5,-34,62,-34</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-34,35.5,-33.5</points>
<intersection>-34 2</intersection>
<intersection>-33.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-33.5,35.5,-33.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-34,42.5,-34</points>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-33.5,16.5,-32</points>
<intersection>-33.5 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-32,16.5,-32</points>
<connection>
<GID>93</GID>
<name>N_in1</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16.5,-33.5,22.5,-33.5</points>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>55,-4</position>
<gparam>LABEL_TEXT RIGHT SHIFT REGISTER (SIPO)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AE_DFF_LOW</type>
<position>28.5,-26</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>58 </output>
<input>
<ID>clock</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>99</ID>
<type>AE_DFF_LOW</type>
<position>45,-26</position>
<input>
<ID>IN_0</ID>58 </input>
<output>
<ID>OUT_0</ID>59 </output>
<input>
<ID>clock</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>101</ID>
<type>AE_DFF_LOW</type>
<position>58.5,-26</position>
<input>
<ID>IN_0</ID>59 </input>
<output>
<ID>OUT_0</ID>60 </output>
<input>
<ID>clock</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>103</ID>
<type>AE_DFF_LOW</type>
<position>73.5,-26</position>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUT_0</ID>61 </output>
<input>
<ID>clock</ID>56 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_TOGGLE</type>
<position>9.5,-18.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>107</ID>
<type>BB_CLOCK</type>
<position>8.5,-32</position>
<output>
<ID>CLK</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>109</ID>
<type>GA_LED</type>
<position>36.5,-12.5</position>
<input>
<ID>N_in2</ID>58 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>GA_LED</type>
<position>51,-12</position>
<input>
<ID>N_in2</ID>59 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>GA_LED</type>
<position>62.5,-12</position>
<input>
<ID>N_in2</ID>60 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>GA_LED</type>
<position>85,-24</position>
<input>
<ID>N_in0</ID>61 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,-32,70.5,-32</points>
<connection>
<GID>107</GID>
<name>CLK</name></connection>
<intersection>25.5 5</intersection>
<intersection>42 4</intersection>
<intersection>55.5 7</intersection>
<intersection>70.5 9</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>42,-32,42,-27</points>
<connection>
<GID>99</GID>
<name>clock</name></connection>
<intersection>-32 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>25.5,-32,25.5,-27</points>
<connection>
<GID>97</GID>
<name>clock</name></connection>
<intersection>-32 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>55.5,-32,55.5,-27</points>
<connection>
<GID>101</GID>
<name>clock</name></connection>
<intersection>-32 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>70.5,-32,70.5,-27</points>
<connection>
<GID>103</GID>
<name>clock</name></connection>
<intersection>-32 1</intersection></vsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-24,18.5,-18.5</points>
<intersection>-24 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-24,25.5,-24</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-18.5,18.5,-18.5</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-24,42,-24</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<connection>
<GID>97</GID>
<name>OUT_0</name></connection>
<intersection>36.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36.5,-24,36.5,-13.5</points>
<connection>
<GID>109</GID>
<name>N_in2</name></connection>
<intersection>-24 1</intersection></vsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-24,55.5,-24</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<intersection>51 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>51,-24,51,-13</points>
<connection>
<GID>111</GID>
<name>N_in2</name></connection>
<intersection>-24 1</intersection></vsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61.5,-24,70.5,-24</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<intersection>62.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>62.5,-24,62.5,-13</points>
<connection>
<GID>113</GID>
<name>N_in2</name></connection>
<intersection>-24 1</intersection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76.5,-24,84,-24</points>
<connection>
<GID>115</GID>
<name>N_in0</name></connection>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection></hsegment></shape></wire></page 6>
<page 7>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>55,-4.5</position>
<gparam>LABEL_TEXT LEFT SHIFT  REGISTER (SIPO)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>AE_DFF_LOW</type>
<position>25,-26</position>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>67 </output>
<input>
<ID>clock</ID>62 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>121</ID>
<type>AE_DFF_LOW</type>
<position>44.5,-26</position>
<input>
<ID>IN_0</ID>65 </input>
<output>
<ID>OUT_0</ID>66 </output>
<input>
<ID>clock</ID>62 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>123</ID>
<type>AE_DFF_LOW</type>
<position>62,-26</position>
<input>
<ID>IN_0</ID>64 </input>
<output>
<ID>OUT_0</ID>65 </output>
<input>
<ID>clock</ID>62 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>125</ID>
<type>AE_DFF_LOW</type>
<position>79,-25.5</position>
<input>
<ID>IN_0</ID>63 </input>
<output>
<ID>OUT_0</ID>64 </output>
<input>
<ID>clock</ID>62 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_TOGGLE</type>
<position>96,-38</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>129</ID>
<type>BB_CLOCK</type>
<position>97,-24</position>
<output>
<ID>CLK</ID>62 </output>
<gparam>angle 180</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>131</ID>
<type>GA_LED</type>
<position>69.5,-41</position>
<input>
<ID>N_in3</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>GA_LED</type>
<position>8.5,-26.5</position>
<input>
<ID>N_in1</ID>67 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>GA_LED</type>
<position>35.5,-40.5</position>
<input>
<ID>N_in3</ID>66 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>GA_LED</type>
<position>56,-41</position>
<input>
<ID>N_in3</ID>65 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87.5,-24,87.5,-13.5</points>
<intersection>-24 2</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-13.5,87.5,-13.5</points>
<intersection>28 8</intersection>
<intersection>47.5 6</intersection>
<intersection>65 3</intersection>
<intersection>82 5</intersection>
<intersection>87.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>87.5,-24,93,-24</points>
<connection>
<GID>129</GID>
<name>CLK</name></connection>
<intersection>87.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>65,-25,65,-13.5</points>
<connection>
<GID>123</GID>
<name>clock</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>82,-24.5,82,-13.5</points>
<connection>
<GID>125</GID>
<name>clock</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>47.5,-25,47.5,-13.5</points>
<connection>
<GID>121</GID>
<name>clock</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>28,-25,28,-13.5</points>
<connection>
<GID>119</GID>
<name>clock</name></connection>
<intersection>-13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-38,88,-27.5</points>
<intersection>-38 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-27.5,88,-27.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>88,-38,94,-38</points>
<connection>
<GID>127</GID>
<name>OUT_0</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-28,70.5,-27.5</points>
<intersection>-28 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65,-28,70.5,-28</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>69.5 3</intersection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-27.5,76,-27.5</points>
<connection>
<GID>125</GID>
<name>OUT_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>69.5,-40,69.5,-28</points>
<connection>
<GID>131</GID>
<name>N_in3</name></connection>
<intersection>-28 1</intersection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>47.5,-28,59,-28</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection>
<intersection>56 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>56,-40,56,-28</points>
<connection>
<GID>137</GID>
<name>N_in3</name></connection>
<intersection>-28 1</intersection></vsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-28,41.5,-28</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<connection>
<GID>121</GID>
<name>OUT_0</name></connection>
<intersection>35.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>35.5,-39.5,35.5,-28</points>
<connection>
<GID>135</GID>
<name>N_in3</name></connection>
<intersection>-28 1</intersection></vsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-28,15.5,-26.5</points>
<intersection>-28 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,-28,22,-28</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-26.5,15.5,-26.5</points>
<connection>
<GID>133</GID>
<name>N_in1</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire></page 7>
<page 8>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>55.5,-4</position>
<gparam>LABEL_TEXT RIGHT SHIFT REGISTER (PIPO)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>AE_DFF_LOW</type>
<position>25,-26</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>73 </output>
<input>
<ID>clock</ID>68 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>143</ID>
<type>AE_DFF_LOW</type>
<position>42.5,-25.5</position>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>74 </output>
<input>
<ID>clock</ID>68 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>145</ID>
<type>AE_DFF_LOW</type>
<position>59,-25.5</position>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>75 </output>
<input>
<ID>clock</ID>68 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>147</ID>
<type>AE_DFF_LOW</type>
<position>75,-26</position>
<input>
<ID>IN_0</ID>72 </input>
<output>
<ID>OUT_0</ID>76 </output>
<input>
<ID>clock</ID>68 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>149</ID>
<type>BB_CLOCK</type>
<position>7,-26.5</position>
<output>
<ID>CLK</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>151</ID>
<type>GA_LED</type>
<position>31.5,-45</position>
<input>
<ID>N_in2</ID>73 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>GA_LED</type>
<position>50,-45.5</position>
<input>
<ID>N_in3</ID>74 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>GA_LED</type>
<position>65,-46</position>
<input>
<ID>N_in3</ID>75 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>GA_LED</type>
<position>80.5,-46.5</position>
<input>
<ID>N_in3</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>AA_TOGGLE</type>
<position>18.5,-12</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_TOGGLE</type>
<position>37,-13</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>163</ID>
<type>AA_TOGGLE</type>
<position>54.5,-11.5</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_TOGGLE</type>
<position>69.5,-12</position>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-35,16.5,-26.5</points>
<intersection>-35 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-35,72,-35</points>
<intersection>16.5 0</intersection>
<intersection>22 4</intersection>
<intersection>39.5 3</intersection>
<intersection>56 6</intersection>
<intersection>72 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-26.5,16.5,-26.5</points>
<connection>
<GID>149</GID>
<name>CLK</name></connection>
<intersection>16.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>39.5,-35,39.5,-26.5</points>
<connection>
<GID>143</GID>
<name>clock</name></connection>
<intersection>-35 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>22,-35,22,-27</points>
<connection>
<GID>141</GID>
<name>clock</name></connection>
<intersection>-35 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>56,-35,56,-26.5</points>
<connection>
<GID>145</GID>
<name>clock</name></connection>
<intersection>-35 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>72,-35,72,-27</points>
<connection>
<GID>147</GID>
<name>clock</name></connection>
<intersection>-35 1</intersection></vsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-24,18.5,-14</points>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18.5,-24,22,-24</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-23.5,37,-15</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37,-23.5,39.5,-23.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>37 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-23.5,54.5,-13.5</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-23.5,56,-23.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-24,69.5,-14</points>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-24,72,-24</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-46,31.5,-24</points>
<connection>
<GID>151</GID>
<name>N_in2</name></connection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-24,31.5,-24</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-44.5,50,-23.5</points>
<connection>
<GID>153</GID>
<name>N_in3</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45.5,-23.5,50,-23.5</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-45,65,-23.5</points>
<connection>
<GID>155</GID>
<name>N_in3</name></connection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-23.5,65,-23.5</points>
<connection>
<GID>145</GID>
<name>OUT_0</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-45.5,80.5,-24</points>
<connection>
<GID>157</GID>
<name>N_in3</name></connection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-24,80.5,-24</points>
<connection>
<GID>147</GID>
<name>OUT_0</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire></page 8>
<page 9>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport>
<gate>
<ID>193</ID>
<type>AA_TOGGLE</type>
<position>44.5,-43.5</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>195</ID>
<type>GA_LED</type>
<position>17.5,-44.5</position>
<input>
<ID>N_in3</ID>87 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>GA_LED</type>
<position>36,-43</position>
<input>
<ID>N_in3</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>167</ID>
<type>AA_LABEL</type>
<position>55.5,-3.5</position>
<gparam>LABEL_TEXT LEFT SHIFT REGISTER (PIPO)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>AE_DFF_LOW</type>
<position>27,-26</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>87 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>171</ID>
<type>AE_DFF_LOW</type>
<position>41.5,-26</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>88 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>173</ID>
<type>AE_DFF_LOW</type>
<position>56.5,-26</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>84 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>175</ID>
<type>AE_DFF_LOW</type>
<position>74.5,-26.5</position>
<input>
<ID>IN_0</ID>78 </input>
<output>
<ID>OUT_0</ID>82 </output>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_TOGGLE</type>
<position>85,-42</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>179</ID>
<type>BB_CLOCK</type>
<position>95,-26</position>
<output>
<ID>CLK</ID>77 </output>
<gparam>angle 180</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_TOGGLE</type>
<position>30,-44.5</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>187</ID>
<type>GA_LED</type>
<position>66.5,-43.5</position>
<input>
<ID>N_in3</ID>82 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>189</ID>
<type>AA_TOGGLE</type>
<position>61,-43.5</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>191</ID>
<type>GA_LED</type>
<position>50,-43</position>
<input>
<ID>N_in3</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-26,84,-11.5</points>
<intersection>-26 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-11.5,84,-11.5</points>
<intersection>30 7</intersection>
<intersection>44.5 8</intersection>
<intersection>59.5 3</intersection>
<intersection>77.5 6</intersection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84,-26,91,-26</points>
<connection>
<GID>179</GID>
<name>CLK</name></connection>
<intersection>84 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>59.5,-25,59.5,-11.5</points>
<connection>
<GID>173</GID>
<name>clock</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>77.5,-25.5,77.5,-11.5</points>
<connection>
<GID>175</GID>
<name>clock</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>30,-25,30,-11.5</points>
<connection>
<GID>169</GID>
<name>clock</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>44.5,-25,44.5,-11.5</points>
<connection>
<GID>171</GID>
<name>clock</name></connection>
<intersection>-11.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-40,85,-28.5</points>
<connection>
<GID>177</GID>
<name>OUT_0</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77.5,-28.5,85,-28.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-42.5,66.5,-28.5</points>
<connection>
<GID>187</GID>
<name>N_in3</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-28.5,71.5,-28.5</points>
<connection>
<GID>175</GID>
<name>OUT_0</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-41.5,61,-28</points>
<connection>
<GID>189</GID>
<name>OUT_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-28,61,-28</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-42,50,-28</points>
<connection>
<GID>191</GID>
<name>N_in3</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-28,53.5,-28</points>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-41.5,44.5,-28</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-42.5,30,-28</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<connection>
<GID>185</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-43.5,17.5,-28</points>
<connection>
<GID>195</GID>
<name>N_in3</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-28,24,-28</points>
<connection>
<GID>169</GID>
<name>OUT_0</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-42,36,-28</points>
<connection>
<GID>197</GID>
<name>N_in3</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-28,38.5,-28</points>
<connection>
<GID>171</GID>
<name>OUT_0</name></connection>
<intersection>36 0</intersection></hsegment></shape></wire></page 9></circuit>