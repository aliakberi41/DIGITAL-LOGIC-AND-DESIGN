<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,3,122.4,-57.5</PageViewport>
<gate>
<ID>2</ID>
<type>BA_DECODER_2x4</type>
<position>36.5,-14</position>
<input>
<ID>ENABLE</ID>1 </input>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT_0</ID>7 </output>
<output>
<ID>OUT_1</ID>6 </output>
<output>
<ID>OUT_2</ID>5 </output>
<output>
<ID>OUT_3</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>13,-4</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>11.5,-11.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>11.5,-17</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>69,-7</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>70.5,-13</position>
<input>
<ID>N_in0</ID>5 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>70.5,-18</position>
<input>
<ID>N_in0</ID>6 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>71,-23.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>34,-30</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_AND2</type>
<position>34,-37.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>34,-45.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>34.5,-54</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>9.5,-27</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>9.5,-35.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_INVERTER</type>
<position>19.5,-27.5</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_INVERTER</type>
<position>19.5,-35.5</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>58.5,-28.5</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>59,-37.5</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>GA_LED</type>
<position>59.5,-45.5</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>GA_LED</type>
<position>60,-54</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>8,-22.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>7.5,-39</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>71.5,-28</position>
<gparam>LABEL_TEXT D0=A'B'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>72,-53.5</position>
<gparam>LABEL_TEXT D3=AB</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_LABEL</type>
<position>71,-36.5</position>
<gparam>LABEL_TEXT D1=A'B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>71.5,-44.5</position>
<gparam>LABEL_TEXT D2=AB'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>54.5,0.5</position>
<gparam>LABEL_TEXT DECODER</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>24.5,-24.5</position>
<gparam>LABEL_TEXT A'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>24.5,-38</position>
<gparam>LABEL_TEXT B'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>101.5,-36</position>
<gparam>LABEL_TEXT (2 TO 4 LINE DECODER)</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-12.5,28,-4</points>
<intersection>-12.5 1</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-12.5,33.5,-12.5</points>
<connection>
<GID>2</GID>
<name>ENABLE</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,-4,28,-4</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-14.5,24,-11.5</points>
<intersection>-14.5 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-14.5,33.5,-14.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-11.5,24,-11.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>24 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-20,27.5,-17</points>
<intersection>-20 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-20,33.5,-20</points>
<intersection>27.5 0</intersection>
<intersection>33.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-17,27.5,-17</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33.5,-20,33.5,-15.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-12.5,43.5,-7</points>
<intersection>-12.5 2</intersection>
<intersection>-7 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-7,68,-7</points>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39.5,-12.5,43.5,-12.5</points>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-13.5,43.5,-13</points>
<intersection>-13.5 2</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-13,69.5,-13</points>
<connection>
<GID>12</GID>
<name>N_in0</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39.5,-13.5,43.5,-13.5</points>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-18,43.5,-14.5</points>
<intersection>-18 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-18,69.5,-18</points>
<connection>
<GID>14</GID>
<name>N_in0</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39.5,-14.5,43.5,-14.5</points>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-23.5,43.5,-15.5</points>
<intersection>-23.5 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-23.5,70,-23.5</points>
<connection>
<GID>16</GID>
<name>N_in0</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39.5,-15.5,43.5,-15.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-30.5,14,-27</points>
<intersection>-30.5 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,-30.5,16.5,-30.5</points>
<intersection>3.5 4</intersection>
<intersection>14 0</intersection>
<intersection>16.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-27,14,-27</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>14 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16.5,-30.5,16.5,-27.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>-30.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>3.5,-44.5,3.5,-30.5</points>
<intersection>-44.5 5</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>3.5,-44.5,31,-44.5</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>3.5 4</intersection>
<intersection>23 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>23,-53,23,-44.5</points>
<intersection>-53 7</intersection>
<intersection>-44.5 5</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>23,-53,31.5,-53</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>23 6</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>7</ID>
<points>29,-55,29,-38.5</points>
<intersection>-55 12</intersection>
<intersection>-38.5 18</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>11.5,-55,31.5,-55</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>11.5 16</intersection>
<intersection>16.5 17</intersection>
<intersection>29 7</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>11.5,-55,11.5,-35.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-55 12</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>16.5,-55,16.5,-35.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>-55 12</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>29,-38.5,31,-38.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>29 7</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-46.5,26.5,-31</points>
<intersection>-46.5 1</intersection>
<intersection>-35.5 2</intersection>
<intersection>-31 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-46.5,31,-46.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-35.5,26.5,-35.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>26.5,-31,31,-31</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-45.5,58.5,-45.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<connection>
<GID>38</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-29,26.5,-27.5</points>
<intersection>-29 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-29,31,-29</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection>
<intersection>31 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-27.5,26.5,-27.5</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>26.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-36.5,31,-29</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-29 1</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-30,40,-28.5</points>
<intersection>-30 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-28.5,57.5,-28.5</points>
<connection>
<GID>34</GID>
<name>N_in0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37,-30,40,-30</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-37.5,58,-37.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<connection>
<GID>36</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-54,59,-54</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<connection>
<GID>40</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-5.67033,1.19597,116.73,-59.3042</PageViewport>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>49.5,-3</position>
<gparam>LABEL_TEXT ENCODER</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_TOGGLE</type>
<position>12.5,-11.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_TOGGLE</type>
<position>12,-20</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_TOGGLE</type>
<position>12.5,-28.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>12.5,-37.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>AE_OR2</type>
<position>46.5,-18.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>86</ID>
<type>AE_OR2</type>
<position>46.5,-29.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>88</ID>
<type>GA_LED</type>
<position>62,-18</position>
<input>
<ID>N_in0</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>GA_LED</type>
<position>62,-30.5</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>7,-10.5</position>
<gparam>LABEL_TEXT I3</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_LABEL</type>
<position>6.5,-19.5</position>
<gparam>LABEL_TEXT I2</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>6.5,-28</position>
<gparam>LABEL_TEXT I1</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>6.5,-36.5</position>
<gparam>LABEL_TEXT I0</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>79.5,-17.5</position>
<gparam>LABEL_TEXT A=I2+I3</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>79.5,-30</position>
<gparam>LABEL_TEXT B=I1+I3</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-20,28.5,-19.5</points>
<intersection>-20 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-19.5,43.5,-19.5</points>
<connection>
<GID>84</GID>
<name>IN_1</name></connection>
<intersection>28.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-20,28.5,-20</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-17.5,29,-11.5</points>
<intersection>-17.5 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-17.5,43.5,-17.5</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection>
<intersection>37.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-11.5,29,-11.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37.5,-28.5,37.5,-17.5</points>
<intersection>-28.5 4</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37.5,-28.5,43.5,-28.5</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>37.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-30.5,29,-28.5</points>
<intersection>-30.5 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-30.5,43.5,-30.5</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14.5,-28.5,29,-28.5</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-18.5,55,-18</points>
<intersection>-18.5 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-18,61,-18</points>
<connection>
<GID>88</GID>
<name>N_in0</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-18.5,55,-18.5</points>
<connection>
<GID>84</GID>
<name>OUT</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-30.5,55,-29.5</points>
<intersection>-30.5 1</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-30.5,61,-30.5</points>
<connection>
<GID>90</GID>
<name>N_in0</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-29.5,55,-29.5</points>
<connection>
<GID>86</GID>
<name>OUT</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-3.86692,1.35556,118.533,-59.1444</PageViewport>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>53.5,-2.5</position>
<gparam>LABEL_TEXT MULTIPLEXERS</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>AA_MUX_2x1</type>
<position>44.5,-22</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>24 </output>
<input>
<ID>SEL_0</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_TOGGLE</type>
<position>24.5,-16</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_TOGGLE</type>
<position>24.5,-24.5</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_TOGGLE</type>
<position>41,-12.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>114</ID>
<type>GA_LED</type>
<position>68,-20.5</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_AND2</type>
<position>27,-33.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_AND2</type>
<position>27.5,-42.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>AE_OR2</type>
<position>51,-37.5</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_TOGGLE</type>
<position>6.5,-29.5</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_TOGGLE</type>
<position>6.5,-39</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_TOGGLE</type>
<position>6.5,-47.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>130</ID>
<type>GA_LED</type>
<position>65,-37</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_INVERTER</type>
<position>16,-48</position>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_LABEL</type>
<position>1,-29.5</position>
<gparam>LABEL_TEXT I1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>AA_LABEL</type>
<position>1.5,-38.5</position>
<gparam>LABEL_TEXT I0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>1.5,-46.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-19.5,44.5,-12.5</points>
<connection>
<GID>106</GID>
<name>SEL_0</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-12.5,44.5,-12.5</points>
<connection>
<GID>112</GID>
<name>OUT_0</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-21,34.5,-16</points>
<intersection>-21 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-21,42.5,-21</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-16,34.5,-16</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-24.5,34.5,-23</points>
<intersection>-24.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-23,42.5,-23</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-24.5,34.5,-24.5</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-22,56.5,-20.5</points>
<intersection>-22 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-20.5,67,-20.5</points>
<connection>
<GID>114</GID>
<name>N_in0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-22,56.5,-22</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59,-37.5,59,-37</points>
<intersection>-37.5 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-37,64,-37</points>
<connection>
<GID>130</GID>
<name>N_in0</name></connection>
<intersection>59 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-37.5,59,-37.5</points>
<connection>
<GID>120</GID>
<name>OUT</name></connection>
<intersection>59 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-36.5,39,-33.5</points>
<intersection>-36.5 1</intersection>
<intersection>-33.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-36.5,48,-36.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-33.5,39,-33.5</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-42.5,39,-38.5</points>
<intersection>-42.5 2</intersection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-38.5,48,-38.5</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-42.5,39,-42.5</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10.5,-47.5,10.5,-43.5</points>
<intersection>-47.5 2</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-43.5,24.5,-43.5</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>10.5 0</intersection>
<intersection>13 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-47.5,10.5,-47.5</points>
<connection>
<GID>128</GID>
<name>OUT_0</name></connection>
<intersection>10.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>13,-48,13,-43.5</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-43.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-41.5,16.5,-29.5</points>
<intersection>-41.5 1</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-41.5,24.5,-41.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>16.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-29.5,16.5,-29.5</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-39,14,-32.5</points>
<intersection>-39 2</intersection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14,-32.5,24,-32.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-39,14,-39</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-48,21.5,-34.5</points>
<intersection>-48 2</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-34.5,24,-34.5</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,-48,21.5,-48</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>21.5 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,7.48321e-007,122.4,-60.5</PageViewport>
<gate>
<ID>5</ID>
<type>AA_TOGGLE</type>
<position>20,-23.5</position>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>94,-3.5</position>
<gparam>LABEL_TEXT (1*2)</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>20,-33.5</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>20.5,-14.5</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_LABEL</type>
<position>55,-3.5</position>
<gparam>LABEL_TEXT DEMULTIPLEXERS</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>GA_LED</type>
<position>73.5,-16.5</position>
<input>
<ID>N_in0</ID>28 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_AND3</type>
<position>60.5,-16</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>35 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>21</ID>
<type>GA_LED</type>
<position>73.5,-26</position>
<input>
<ID>N_in0</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_AND3</type>
<position>60.5,-31.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>37 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_LABEL</type>
<position>56,-45.5</position>
<gparam>LABEL_TEXT (BY USING ENABLE)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>16.5,-14</position>
<gparam>LABEL_TEXT I</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>15.5,-23</position>
<gparam>LABEL_TEXT E</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>15,-33.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>AA_INVERTER</type>
<position>33,-33.5</position>
<input>
<ID>IN_0</ID>37 </input>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>87,-15.5</position>
<gparam>LABEL_TEXT D0=IES'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>87,-26</position>
<gparam>LABEL_TEXT D1=IES</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-16.5,68,-16</points>
<intersection>-16.5 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-16.5,72.5,-16.5</points>
<connection>
<GID>17</GID>
<name>N_in0</name></connection>
<intersection>68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-16,68,-16</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-31.5,68,-26</points>
<intersection>-31.5 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-26,72.5,-26</points>
<connection>
<GID>21</GID>
<name>N_in0</name></connection>
<intersection>68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-31.5,68,-31.5</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-14.5,40,-14</points>
<intersection>-14.5 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-14,57.5,-14</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>40 0</intersection>
<intersection>53 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-14.5,40,-14.5</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>40 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>53,-29.5,53,-14</points>
<intersection>-29.5 4</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>53,-29.5,57.5,-29.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>53 3</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-33.5,46.5,-18</points>
<intersection>-33.5 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-18,57.5,-18</points>
<connection>
<GID>19</GID>
<name>IN_2</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36,-33.5,46.5,-33.5</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-38.5,57.5,-38.5</points>
<intersection>22 6</intersection>
<intersection>30 5</intersection>
<intersection>57.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>57.5,-38.5,57.5,-33.5</points>
<connection>
<GID>25</GID>
<name>IN_2</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>30,-38.5,30,-33.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>22,-38.5,22,-33.5</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<intersection>-38.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-23.5,39.5,-16</points>
<intersection>-23.5 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-16,57.5,-16</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection>
<intersection>53 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-23.5,39.5,-23.5</points>
<connection>
<GID>5</GID>
<name>OUT_0</name></connection>
<intersection>39.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>53,-31.5,53,-16</points>
<intersection>-31.5 4</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>53,-31.5,57.5,-31.5</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>53 3</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-13.0999,2.74917,109.3,-57.7508</PageViewport>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>44.5,0</position>
<gparam>LABEL_TEXT DECODERS</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>76,-8.5</position>
<input>
<ID>N_in0</ID>60 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>GA_LED</type>
<position>76,-16</position>
<input>
<ID>N_in0</ID>61 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>76,-22.5</position>
<input>
<ID>N_in0</ID>62 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>GA_LED</type>
<position>76,-29</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>GA_LED</type>
<position>76,-34</position>
<input>
<ID>N_in0</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>GA_LED</type>
<position>76,-40</position>
<input>
<ID>N_in0</ID>65 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>242</ID>
<type>AA_LABEL</type>
<position>87,-8</position>
<gparam>LABEL_TEXT D0=X'Y'Z'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>GA_LED</type>
<position>76,-46.5</position>
<input>
<ID>N_in0</ID>66 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>244</ID>
<type>AA_LABEL</type>
<position>87,-15</position>
<gparam>LABEL_TEXT D1=X'Y'Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>246</ID>
<type>AA_LABEL</type>
<position>87.5,-22</position>
<gparam>LABEL_TEXT D2=X'YZ'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>GA_LED</type>
<position>76,-53.5</position>
<input>
<ID>N_in0</ID>67 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>248</ID>
<type>AA_LABEL</type>
<position>88,-28.5</position>
<gparam>LABEL_TEXT D3=X'YZ</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>250</ID>
<type>AA_LABEL</type>
<position>88,-33.5</position>
<gparam>LABEL_TEXT D4=XY'Z'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>252</ID>
<type>AA_LABEL</type>
<position>88,-39</position>
<gparam>LABEL_TEXT D5=XY'Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>254</ID>
<type>AA_LABEL</type>
<position>88.5,-45.5</position>
<gparam>LABEL_TEXT D6=XYZ'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>256</ID>
<type>AA_LABEL</type>
<position>88.5,-53</position>
<gparam>LABEL_TEXT D7=XYZ</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>0.5,-7.5</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>258</ID>
<type>AA_LABEL</type>
<position>-3.5,-7</position>
<gparam>LABEL_TEXT E</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_TOGGLE</type>
<position>1.5,-15.5</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>260</ID>
<type>AA_LABEL</type>
<position>-4.5,-15</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>262</ID>
<type>AA_LABEL</type>
<position>-4,-26.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_TOGGLE</type>
<position>1.5,-27</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>264</ID>
<type>AA_LABEL</type>
<position>-4,-37</position>
<gparam>LABEL_TEXT Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>BE_DECODER_3x8</type>
<position>46,-14.5</position>
<input>
<ID>ENABLE</ID>68 </input>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>70 </input>
<input>
<ID>IN_2</ID>69 </input>
<output>
<ID>OUT_0</ID>67 </output>
<output>
<ID>OUT_1</ID>66 </output>
<output>
<ID>OUT_2</ID>65 </output>
<output>
<ID>OUT_3</ID>64 </output>
<output>
<ID>OUT_4</ID>63 </output>
<output>
<ID>OUT_5</ID>62 </output>
<output>
<ID>OUT_6</ID>61 </output>
<output>
<ID>OUT_7</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>119</ID>
<type>AA_TOGGLE</type>
<position>1.5,-37.5</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>12.5,-46.5</position>
<gparam>LABEL_TEXT 3*8 LINE DECODER</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-11,62,-6</points>
<intersection>-11 2</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62,-6,75,-6</points>
<intersection>62 0</intersection>
<intersection>75 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-11,62,-11</points>
<connection>
<GID>115</GID>
<name>OUT_7</name></connection>
<intersection>62 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75,-8.5,75,-6</points>
<connection>
<GID>27</GID>
<name>N_in0</name></connection>
<intersection>-6 1</intersection></vsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-20,63,-12</points>
<intersection>-20 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-20,75,-20</points>
<intersection>63 0</intersection>
<intersection>75 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-12,63,-12</points>
<connection>
<GID>115</GID>
<name>OUT_6</name></connection>
<intersection>63 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>75,-20,75,-16</points>
<connection>
<GID>31</GID>
<name>N_in0</name></connection>
<intersection>-20 1</intersection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-22.5,61,-13</points>
<intersection>-22.5 1</intersection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-22.5,75,-22.5</points>
<connection>
<GID>35</GID>
<name>N_in0</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-13,61,-13</points>
<connection>
<GID>115</GID>
<name>OUT_5</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-29,59.5,-14</points>
<intersection>-29 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-29,75,-29</points>
<connection>
<GID>39</GID>
<name>N_in0</name></connection>
<intersection>59.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-14,59.5,-14</points>
<connection>
<GID>115</GID>
<name>OUT_4</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58,-34,58,-15</points>
<intersection>-34 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-34,75,-34</points>
<connection>
<GID>43</GID>
<name>N_in0</name></connection>
<intersection>58 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-15,58,-15</points>
<connection>
<GID>115</GID>
<name>OUT_3</name></connection>
<intersection>58 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57,-40,57,-16</points>
<intersection>-40 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>57,-40,75,-40</points>
<connection>
<GID>47</GID>
<name>N_in0</name></connection>
<intersection>57 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-16,57,-16</points>
<connection>
<GID>115</GID>
<name>OUT_2</name></connection>
<intersection>57 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-46.5,56,-17</points>
<intersection>-46.5 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-46.5,75,-46.5</points>
<connection>
<GID>51</GID>
<name>N_in0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-17,56,-17</points>
<connection>
<GID>115</GID>
<name>OUT_1</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-49,54,-18</points>
<intersection>-49 1</intersection>
<intersection>-18 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-49,72.5,-49</points>
<intersection>54 0</intersection>
<intersection>72.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49,-18,54,-18</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>54 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>72.5,-53.5,72.5,-49</points>
<intersection>-53.5 4</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>72.5,-53.5,75,-53.5</points>
<connection>
<GID>55</GID>
<name>N_in0</name></connection>
<intersection>72.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-11,27,-7.5</points>
<intersection>-11 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-11,43,-11</points>
<connection>
<GID>115</GID>
<name>ENABLE</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>2.5,-7.5,27,-7.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3.5,-15.5,43,-15.5</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>43 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43,-16,43,-15.5</points>
<connection>
<GID>115</GID>
<name>IN_2</name></connection>
<intersection>-15.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-27,27,-17</points>
<intersection>-27 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,-17,43,-17</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>27 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-27,27,-27</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>27 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-37.5,32.5,-18</points>
<intersection>-37.5 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-18,43,-18</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-37.5,32.5,-37.5</points>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>0.342031,-0.539213,122.742,-61.0392</PageViewport>
<gate>
<ID>194</ID>
<type>AA_LABEL</type>
<position>91.5,-11</position>
<gparam>LABEL_TEXT D1=X'Y'Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>196</ID>
<type>AA_LABEL</type>
<position>92,-19</position>
<gparam>LABEL_TEXT D2=X'YZ'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>198</ID>
<type>AA_LABEL</type>
<position>91.5,-26.5</position>
<gparam>LABEL_TEXT D3=X'YZ</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>200</ID>
<type>AA_LABEL</type>
<position>92.5,-34</position>
<gparam>LABEL_TEXT D4=XY'Z'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>AA_LABEL</type>
<position>92.5,-42</position>
<gparam>LABEL_TEXT D5=XY'Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>204</ID>
<type>AA_LABEL</type>
<position>93,-48.5</position>
<gparam>LABEL_TEXT D6=XYZ'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>206</ID>
<type>AA_LABEL</type>
<position>92.5,-56</position>
<gparam>LABEL_TEXT D7=XYZ</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>AA_LABEL</type>
<position>19,-53.5</position>
<gparam>LABEL_TEXT 3*8 LINE DECODER</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>AA_AND3</type>
<position>65,-4.5</position>
<input>
<ID>IN_0</ID>87 </input>
<input>
<ID>IN_1</ID>86 </input>
<input>
<ID>IN_2</ID>88 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>137</ID>
<type>AA_AND3</type>
<position>65,-12.5</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>86 </input>
<input>
<ID>IN_2</ID>80 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_AND3</type>
<position>65,-20</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>81 </input>
<input>
<ID>IN_2</ID>87 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_AND3</type>
<position>65,-27.5</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>81 </input>
<input>
<ID>IN_2</ID>80 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_AND3</type>
<position>65,-35</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>86 </input>
<input>
<ID>IN_2</ID>87 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>146</ID>
<type>AA_AND3</type>
<position>65,-43</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>86 </input>
<input>
<ID>IN_2</ID>80 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_AND3</type>
<position>65,-50</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>81 </input>
<input>
<ID>IN_2</ID>87 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_AND3</type>
<position>65,-57</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>81 </input>
<input>
<ID>IN_2</ID>80 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>152</ID>
<type>GA_LED</type>
<position>79,-4.5</position>
<input>
<ID>N_in0</ID>79 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>79,-11.5</position>
<input>
<ID>N_in0</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>GA_LED</type>
<position>79.5,-20</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>GA_LED</type>
<position>79.5,-27</position>
<input>
<ID>N_in0</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>GA_LED</type>
<position>79.5,-34.5</position>
<input>
<ID>N_in0</ID>75 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>GA_LED</type>
<position>79.5,-42</position>
<input>
<ID>N_in0</ID>74 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>GA_LED</type>
<position>79.5,-48.5</position>
<input>
<ID>N_in0</ID>73 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>GA_LED</type>
<position>79.5,-57</position>
<input>
<ID>N_in0</ID>72 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AA_TOGGLE</type>
<position>11,-12.5</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_TOGGLE</type>
<position>11,-28</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_TOGGLE</type>
<position>11,-44.5</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>174</ID>
<type>AA_INVERTER</type>
<position>21.5,-12.5</position>
<input>
<ID>IN_0</ID>80 </input>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_INVERTER</type>
<position>22.5,-28</position>
<input>
<ID>IN_0</ID>81 </input>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_INVERTER</type>
<position>23,-44.5</position>
<input>
<ID>IN_0</ID>82 </input>
<output>
<ID>OUT_0</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>91.5,-4</position>
<gparam>LABEL_TEXT D0=X'Y'Z'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>AA_LABEL</type>
<position>6.5,-43.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>6,-27.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>21.5,-16.5</position>
<gparam>LABEL_TEXT Z'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>188</ID>
<type>AA_LABEL</type>
<position>23,-48.5</position>
<gparam>LABEL_TEXT X'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>AA_LABEL</type>
<position>22,-32.5</position>
<gparam>LABEL_TEXT Y'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>192</ID>
<type>AA_LABEL</type>
<position>6.5,-12</position>
<gparam>LABEL_TEXT Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-57,78.5,-57</points>
<connection>
<GID>166</GID>
<name>N_in0</name></connection>
<connection>
<GID>150</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-50,73,-48.5</points>
<intersection>-50 2</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-48.5,78.5,-48.5</points>
<connection>
<GID>164</GID>
<name>N_in0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-50,73,-50</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-43,73,-42</points>
<intersection>-43 2</intersection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-42,78.5,-42</points>
<connection>
<GID>162</GID>
<name>N_in0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-43,73,-43</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-35,73,-34.5</points>
<intersection>-35 2</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-34.5,78.5,-34.5</points>
<connection>
<GID>160</GID>
<name>N_in0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-35,73,-35</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-27.5,73,-27</points>
<intersection>-27.5 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-27,78.5,-27</points>
<connection>
<GID>158</GID>
<name>N_in0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-27.5,73,-27.5</points>
<connection>
<GID>142</GID>
<name>OUT</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-20,78.5,-20</points>
<connection>
<GID>156</GID>
<name>N_in0</name></connection>
<connection>
<GID>140</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-12.5,73,-11.5</points>
<intersection>-12.5 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-11.5,78,-11.5</points>
<connection>
<GID>154</GID>
<name>N_in0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-12.5,73,-12.5</points>
<connection>
<GID>137</GID>
<name>OUT</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-4.5,78,-4.5</points>
<connection>
<GID>152</GID>
<name>N_in0</name></connection>
<connection>
<GID>133</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-15,62,-15</points>
<intersection>13 3</intersection>
<intersection>18.5 4</intersection>
<intersection>42 2</intersection>
<intersection>62 8</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>42,-45,42,-15</points>
<intersection>-45 10</intersection>
<intersection>-29.5 7</intersection>
<intersection>-15 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>13,-15,13,-12.5</points>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection>
<intersection>-15 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>18.5,-15,18.5,-12.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>42,-29.5,62,-29.5</points>
<connection>
<GID>142</GID>
<name>IN_2</name></connection>
<intersection>42 2</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>62,-15,62,-14.5</points>
<connection>
<GID>137</GID>
<name>IN_2</name></connection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>37.5,-45,62,-45</points>
<connection>
<GID>146</GID>
<name>IN_2</name></connection>
<intersection>37.5 11</intersection>
<intersection>42 2</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>37.5,-59,37.5,-45</points>
<intersection>-59 12</intersection>
<intersection>-45 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>37.5,-59,62,-59</points>
<connection>
<GID>150</GID>
<name>IN_2</name></connection>
<intersection>37.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-20,62,-20</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<intersection>13 5</intersection>
<intersection>19.5 4</intersection>
<intersection>47 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>19.5,-28,19.5,-20</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>-20 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>13,-28,13,-20</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<intersection>-20 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>47,-50,47,-20</points>
<intersection>-50 9</intersection>
<intersection>-27.5 7</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>47,-27.5,62,-27.5</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>47 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>42,-50,62,-50</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<intersection>42 10</intersection>
<intersection>47 6</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>42,-57,42,-50</points>
<intersection>-57 11</intersection>
<intersection>-50 9</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>42,-57,62,-57</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>42 10</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-35,36,-35</points>
<intersection>13 6</intersection>
<intersection>20 5</intersection>
<intersection>36 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-35,36,-33</points>
<intersection>-35 1</intersection>
<intersection>-33 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36,-33,62,-33</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>36 3</intersection>
<intersection>47 7</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>20,-44.5,20,-35</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>13,-44.5,13,-35</points>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<intersection>-35 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>47,-41,47,-33</points>
<intersection>-41 8</intersection>
<intersection>-33 4</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>42,-41,62,-41</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>42 9</intersection>
<intersection>47 7</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>42,-48,42,-41</points>
<intersection>-48 10</intersection>
<intersection>-41 8</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>42,-48,62,-48</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>42 9</intersection>
<intersection>47 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>47,-55,47,-48</points>
<intersection>-55 12</intersection>
<intersection>-48 10</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>47,-55,62,-55</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>47 11</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-28,31,-4.5</points>
<intersection>-28 2</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-4.5,62,-4.5</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>31 0</intersection>
<intersection>53 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25.5,-28,31,-28</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<intersection>31 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>53,-12.5,53,-4.5</points>
<intersection>-12.5 4</intersection>
<intersection>-4.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-12.5,62,-12.5</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<intersection>50.5 5</intersection>
<intersection>53 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>50.5,-35,50.5,-12.5</points>
<intersection>-35 6</intersection>
<intersection>-12.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>50.5,-35,62,-35</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>50.5 5</intersection>
<intersection>57 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>57,-43,57,-35</points>
<intersection>-43 8</intersection>
<intersection>-35 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>57,-43,62,-43</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>57 7</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-12.5,29.5,-2.5</points>
<intersection>-12.5 1</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-12.5,29.5,-12.5</points>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-2.5,62,-2.5</points>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>29.5 0</intersection>
<intersection>50.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50.5,-52,50.5,-2.5</points>
<intersection>-52 8</intersection>
<intersection>-37 6</intersection>
<intersection>-22 4</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-22,62,-22</points>
<connection>
<GID>140</GID>
<name>IN_2</name></connection>
<intersection>50.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>50.5,-37,62,-37</points>
<connection>
<GID>144</GID>
<name>IN_2</name></connection>
<intersection>50.5 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>50.5,-52,62,-52</points>
<connection>
<GID>148</GID>
<name>IN_2</name></connection>
<intersection>50.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-44.5,32.5,-6.5</points>
<intersection>-44.5 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-6.5,62,-6.5</points>
<connection>
<GID>133</GID>
<name>IN_2</name></connection>
<intersection>32.5 0</intersection>
<intersection>56 3</intersection>
<intersection>60.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-44.5,32.5,-44.5</points>
<connection>
<GID>178</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>56,-25.5,56,-6.5</points>
<intersection>-25.5 6</intersection>
<intersection>-18 4</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>56,-18,62,-18</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>56 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>56,-25.5,62,-25.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>56 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>60.5,-10.5,60.5,-6.5</points>
<intersection>-10.5 8</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>60.5,-10.5,62,-10.5</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<intersection>60.5 7</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>8.88178e-016,7.48321e-007,122.4,-60.5</PageViewport>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>50.5,-3.5</position>
<gparam>LABEL_TEXT ENCODER</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_TOGGLE</type>
<position>11,-11.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>78,-3.5</position>
<gparam>LABEL_TEXT (8*3)</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>11,-17</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_TOGGLE</type>
<position>11,-23</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_TOGGLE</type>
<position>11,-28.5</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>11,-34.5</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_TOGGLE</type>
<position>11,-39.5</position>
<output>
<ID>OUT_0</ID>42 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>11.5,-44.5</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>11.5,-49</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>79</ID>
<type>AE_OR4</type>
<position>59,-15.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>42 </input>
<input>
<ID>IN_2</ID>43 </input>
<input>
<ID>IN_3</ID>44 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>83</ID>
<type>AE_OR4</type>
<position>59.5,-29</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<input>
<ID>IN_2</ID>43 </input>
<input>
<ID>IN_3</ID>44 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>87</ID>
<type>AA_AND4</type>
<position>-52.5,-28.5</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_OR4</type>
<position>59.5,-43</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>46 </input>
<input>
<ID>IN_2</ID>42 </input>
<input>
<ID>IN_3</ID>44 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>95</ID>
<type>GA_LED</type>
<position>70.5,-15</position>
<input>
<ID>N_in0</ID>36 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>GA_LED</type>
<position>70.5,-28.5</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>GA_LED</type>
<position>70.5,-43.5</position>
<input>
<ID>N_in0</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>6,-11</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>AA_LABEL</type>
<position>6,-17</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>6,-22.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>AA_LABEL</type>
<position>6.5,-28</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>6,-34</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>AA_LABEL</type>
<position>6,-39</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>6.5,-44</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>AA_LABEL</type>
<position>6.5,-48.5</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>147</ID>
<type>AA_LABEL</type>
<position>89,-14</position>
<gparam>LABEL_TEXT X=D4+D5+D6+D7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>AA_LABEL</type>
<position>90,-27.5</position>
<gparam>LABEL_TEXT Y=D2+D3+D6+D7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>AA_LABEL</type>
<position>90.5,-42.5</position>
<gparam>LABEL_TEXT Z=D1+D3+D5+D7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-15.5,66,-15</points>
<intersection>-15.5 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66,-15,69.5,-15</points>
<connection>
<GID>95</GID>
<name>N_in0</name></connection>
<intersection>66 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-15.5,66,-15.5</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<intersection>66 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-29,66.5,-28.5</points>
<intersection>-29 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-28.5,69.5,-28.5</points>
<connection>
<GID>99</GID>
<name>N_in0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-29,66.5,-29</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-43.5,66.5,-43</points>
<intersection>-43.5 1</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-43.5,69.5,-43.5</points>
<connection>
<GID>103</GID>
<name>N_in0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-43,66.5,-43</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-34.5,20,-12.5</points>
<intersection>-34.5 2</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-12.5,56,-12.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-34.5,20,-34.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>20 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>21.5,-39.5,21.5,-14.5</points>
<intersection>-39.5 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-14.5,56,-14.5</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>21.5 0</intersection>
<intersection>37.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-39.5,21.5,-39.5</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>21.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37.5,-44,37.5,-14.5</points>
<intersection>-44 4</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37.5,-44,56.5,-44</points>
<connection>
<GID>91</GID>
<name>IN_2</name></connection>
<intersection>37.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-44.5,23,-16.5</points>
<intersection>-44.5 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-16.5,56,-16.5</points>
<connection>
<GID>79</GID>
<name>IN_2</name></connection>
<intersection>23 0</intersection>
<intersection>50 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-44.5,23,-44.5</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>23 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50,-30,50,-16.5</points>
<intersection>-30 4</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>50,-30,56.5,-30</points>
<connection>
<GID>83</GID>
<name>IN_2</name></connection>
<intersection>50 3</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-49,24.5,-18.5</points>
<intersection>-49 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-18.5,56,-18.5</points>
<connection>
<GID>79</GID>
<name>IN_3</name></connection>
<intersection>24.5 0</intersection>
<intersection>44 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13.5,-49,24.5,-49</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>24.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>44,-32,44,-18.5</points>
<intersection>-32 4</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>44,-32,56.5,-32</points>
<connection>
<GID>83</GID>
<name>IN_3</name></connection>
<intersection>44 3</intersection>
<intersection>50 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>50,-46,50,-32</points>
<intersection>-46 6</intersection>
<intersection>-32 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>50,-46,56.5,-46</points>
<connection>
<GID>91</GID>
<name>IN_3</name></connection>
<intersection>50 5</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-26,34.5,-23</points>
<intersection>-26 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-26,56.5,-26</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-23,34.5,-23</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-28,56.5,-28</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>13 3</intersection>
<intersection>40 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13,-28.5,13,-28</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>-28 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>40,-42,40,-28</points>
<intersection>-42 5</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>40,-42,56.5,-42</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>40 4</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-40,34.5,-17.5</points>
<intersection>-40 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-40,56.5,-40</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-17.5,34.5,-17.5</points>
<intersection>13 3</intersection>
<intersection>34.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13,-17.5,13,-17</points>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection>
<intersection>-17.5 2</intersection></vsegment></shape></wire></page 6>
<page 7>
<PageViewport>0,7.48321e-007,122.4,-60.5</PageViewport>
<gate>
<ID>195</ID>
<type>AA_INVERTER</type>
<position>26.5,-17</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>199</ID>
<type>AA_INVERTER</type>
<position>27,-31</position>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>203</ID>
<type>AA_LABEL</type>
<position>11.5,-16.5</position>
<gparam>LABEL_TEXT I1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>207</ID>
<type>AA_LABEL</type>
<position>12,-30.5</position>
<gparam>LABEL_TEXT I0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>16,-36.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>16,-41</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_TOGGLE</type>
<position>16,-46.5</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>16,-51</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>10,-36</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>10,-40.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>10,-46</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>10,-50.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>AA_LABEL</type>
<position>102.5,-32</position>
<gparam>LABEL_TEXT X=I0'.I1'.D0+</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>104,-36</position>
<gparam>LABEL_TEXT I0.I1'D1+</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>AA_LABEL</type>
<position>105,-40</position>
<gparam>LABEL_TEXT I0'.I1.D2+</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>AA_LABEL</type>
<position>104,-44</position>
<gparam>LABEL_TEXT I0.I1.D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>153</ID>
<type>AA_LABEL</type>
<position>61,-21</position>
<gparam>LABEL_TEXT I0'.I1'.D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>159</ID>
<type>AA_LABEL</type>
<position>59,-3.5</position>
<gparam>LABEL_TEXT MULTIPLEXERS (4*1)</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>60.5,-33</position>
<gparam>LABEL_TEXT I0.I1'D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>AA_TOGGLE</type>
<position>16,-17</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_TOGGLE</type>
<position>16,-31</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_LABEL</type>
<position>61,-44</position>
<gparam>LABEL_TEXT I0'.I1.D2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>AA_AND3</type>
<position>58,-16</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<input>
<ID>IN_2</ID>57 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_AND3</type>
<position>58.5,-28</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>58 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_LABEL</type>
<position>62,-54.5</position>
<gparam>LABEL_TEXT I0.I1.D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>179</ID>
<type>AA_AND3</type>
<position>58.5,-39</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>59 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>183</ID>
<type>AA_AND3</type>
<position>58.5,-49.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>49 </input>
<input>
<ID>IN_2</ID>83 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>187</ID>
<type>AE_OR4</type>
<position>86,-27</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>54 </input>
<input>
<ID>IN_2</ID>55 </input>
<input>
<ID>IN_3</ID>56 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>191</ID>
<type>GA_LED</type>
<position>98,-27</position>
<input>
<ID>N_in0</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,-27,97,-27</points>
<connection>
<GID>191</GID>
<name>N_in0</name></connection>
<connection>
<GID>187</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-22.5,48,-22.5</points>
<intersection>18 6</intersection>
<intersection>23.5 5</intersection>
<intersection>48 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48,-49.5,48,-22.5</points>
<intersection>-49.5 8</intersection>
<intersection>-37 4</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>48,-37,55.5,-37</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>48 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>23.5,-22.5,23.5,-17</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>-22.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>18,-22.5,18,-17</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>48,-49.5,55.5,-49.5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>48 3</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-31,50.5,-31</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<connection>
<GID>167</GID>
<name>OUT_0</name></connection>
<intersection>44.5 5</intersection>
<intersection>50.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50.5,-31,50.5,-28</points>
<intersection>-31 1</intersection>
<intersection>-28 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-28,55.5,-28</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>50.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>44.5,-39,44.5,-31</points>
<intersection>-39 6</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>44.5,-39,55.5,-39</points>
<connection>
<GID>179</GID>
<name>IN_1</name></connection>
<intersection>44.5 5</intersection>
<intersection>51 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>51,-47.5,51,-39</points>
<intersection>-47.5 8</intersection>
<intersection>-39 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>51,-47.5,55.5,-47.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>51 7</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-17,31.5,-14</points>
<intersection>-17 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-14,55,-14</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>31.5 0</intersection>
<intersection>50.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-17,31.5,-17</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50.5,-26,50.5,-14</points>
<intersection>-26 4</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-26,55.5,-26</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>50.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-31,32.5,-16</points>
<intersection>-31 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-16,55,-16</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30,-31,32.5,-31</points>
<connection>
<GID>199</GID>
<name>OUT_0</name></connection>
<intersection>32.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-24,72,-16</points>
<intersection>-24 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-24,83,-24</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61,-16,72,-16</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-28,72,-26</points>
<intersection>-28 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-26,83,-26</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,-28,72,-28</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-39,73,-28</points>
<intersection>-39 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-28,83,-28</points>
<connection>
<GID>187</GID>
<name>IN_2</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,-39,73,-39</points>
<connection>
<GID>179</GID>
<name>OUT</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-49.5,76,-30</points>
<intersection>-49.5 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-30,83,-30</points>
<connection>
<GID>187</GID>
<name>IN_3</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61.5,-49.5,76,-49.5</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-36.5,36.5,-18</points>
<intersection>-36.5 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-18,55,-18</points>
<connection>
<GID>171</GID>
<name>IN_2</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-36.5,36.5,-36.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-41,39,-30</points>
<intersection>-41 2</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-30,55.5,-30</points>
<connection>
<GID>175</GID>
<name>IN_2</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-41,39,-41</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-46.5,41.5,-41</points>
<intersection>-46.5 2</intersection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-41,55.5,-41</points>
<connection>
<GID>179</GID>
<name>IN_2</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-46.5,41.5,-46.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18,-51,55.5,-51</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>55.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>55.5,-51.5,55.5,-51</points>
<connection>
<GID>183</GID>
<name>IN_2</name></connection>
<intersection>-51 1</intersection></vsegment></shape></wire></page 7>
<page 8>
<PageViewport>-6,6,116.4,-54.5</PageViewport>
<gate>
<ID>193</ID>
<type>AE_MUX_4x1</type>
<position>65,-24.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>89 </input>
<input>
<ID>IN_2</ID>85 </input>
<input>
<ID>IN_3</ID>84 </input>
<output>
<ID>OUT</ID>91 </output>
<input>
<ID>SEL_0</ID>93 </input>
<input>
<ID>SEL_1</ID>92 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_TOGGLE</type>
<position>26.5,-15</position>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_TOGGLE</type>
<position>24,-22.5</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_TOGGLE</type>
<position>25,-29</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_TOGGLE</type>
<position>26.5,-35.5</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>216</ID>
<type>GA_LED</type>
<position>86.5,-23.5</position>
<input>
<ID>N_in0</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>AA_TOGGLE</type>
<position>56,-12.5</position>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_TOGGLE</type>
<position>61,-10.5</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>17.5,-14.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>224</ID>
<type>AA_LABEL</type>
<position>17.5,-22</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>226</ID>
<type>AA_LABEL</type>
<position>18,-28.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>228</ID>
<type>AA_LABEL</type>
<position>18,-35.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>230</ID>
<type>AA_LABEL</type>
<position>54,-9</position>
<gparam>LABEL_TEXT I0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>232</ID>
<type>AA_LABEL</type>
<position>61,-6.5</position>
<gparam>LABEL_TEXT I1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>234</ID>
<type>AA_LABEL</type>
<position>86,-27.5</position>
<gparam>LABEL_TEXT X=I0'.I1'.D0+</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>236</ID>
<type>AA_LABEL</type>
<position>87,-31.5</position>
<gparam>LABEL_TEXT I0.I1'D1+</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>238</ID>
<type>AA_LABEL</type>
<position>88,-36</position>
<gparam>LABEL_TEXT I0'.I1.D2+</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>240</ID>
<type>AA_LABEL</type>
<position>87,-40.5</position>
<gparam>LABEL_TEXT I0.I1.D3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>AA_LABEL</type>
<position>56.5,2</position>
<gparam>LABEL_TEXT MULTIPLEXERS (4*1)</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-21.5,40,-15</points>
<intersection>-21.5 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-21.5,62,-21.5</points>
<connection>
<GID>193</GID>
<name>IN_3</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-15,40,-15</points>
<connection>
<GID>201</GID>
<name>OUT_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-23.5,62,-23.5</points>
<connection>
<GID>193</GID>
<name>IN_2</name></connection>
<intersection>28.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>28.5,-23.5,28.5,-22.5</points>
<intersection>-23.5 1</intersection>
<intersection>-22.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>26,-22.5,28.5,-22.5</points>
<connection>
<GID>209</GID>
<name>OUT_0</name></connection>
<intersection>28.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-29,40,-25.5</points>
<intersection>-29 2</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-25.5,62,-25.5</points>
<connection>
<GID>193</GID>
<name>IN_1</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-29,40,-29</points>
<connection>
<GID>212</GID>
<name>OUT_0</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-35.5,42,-27.5</points>
<intersection>-35.5 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-27.5,62,-27.5</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>42 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-35.5,42,-35.5</points>
<connection>
<GID>214</GID>
<name>OUT_0</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76,-24.5,76,-23.5</points>
<intersection>-24.5 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>76,-23.5,85.5,-23.5</points>
<connection>
<GID>216</GID>
<name>N_in0</name></connection>
<intersection>76 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-24.5,76,-24.5</points>
<connection>
<GID>193</GID>
<name>OUT</name></connection>
<intersection>76 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65,-19.5,65,-12.5</points>
<connection>
<GID>193</GID>
<name>SEL_1</name></connection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58,-12.5,65,-12.5</points>
<connection>
<GID>218</GID>
<name>OUT_0</name></connection>
<intersection>65 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-19.5,66,-10.5</points>
<connection>
<GID>193</GID>
<name>SEL_0</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-10.5,66,-10.5</points>
<connection>
<GID>220</GID>
<name>OUT_0</name></connection>
<intersection>66 0</intersection></hsegment></shape></wire></page 8>
<page 9>
<PageViewport>0,7.48321e-007,122.4,-60.5</PageViewport>
<gate>
<ID>205</ID>
<type>AA_LABEL</type>
<position>13,-29</position>
<gparam>LABEL_TEXT I</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>213</ID>
<type>AA_LABEL</type>
<position>87.5,-18</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>217</ID>
<type>AA_LABEL</type>
<position>88,-29.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>59.5,-4.5</position>
<gparam>LABEL_TEXT DEMULTIPLEXERS(1*2)</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_TOGGLE</type>
<position>17.5,-17</position>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_TOGGLE</type>
<position>16.5,-30.5</position>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_INVERTER</type>
<position>33.5,-17</position>
<input>
<ID>IN_0</ID>94 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>121</ID>
<type>GA_LED</type>
<position>79,-19</position>
<input>
<ID>N_in0</ID>97 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>GA_LED</type>
<position>79,-30</position>
<input>
<ID>N_in0</ID>98 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>AA_AND2</type>
<position>67.5,-18.5</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_AND2</type>
<position>68,-29.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_LABEL</type>
<position>13,-16.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>94</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-17,30.5,-17</points>
<connection>
<GID>72</GID>
<name>OUT_0</name></connection>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>27.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>27.5,-28.5,27.5,-17</points>
<intersection>-28.5 5</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>27.5,-28.5,65,-28.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>27.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-17.5,50.5,-17</points>
<intersection>-17.5 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-17.5,64.5,-17.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-17,50.5,-17</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-30.5,42,-19.5</points>
<intersection>-30.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-19.5,64.5,-19.5</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>42 0</intersection>
<intersection>63.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-30.5,42,-30.5</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<intersection>42 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>63.5,-30.5,63.5,-19.5</points>
<intersection>-30.5 4</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>63.5,-30.5,65,-30.5</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>63.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-19,74,-18.5</points>
<intersection>-19 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-19,78,-19</points>
<connection>
<GID>121</GID>
<name>N_in0</name></connection>
<intersection>74 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-18.5,74,-18.5</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-30,74.5,-29.5</points>
<intersection>-30 1</intersection>
<intersection>-29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-30,78,-30</points>
<connection>
<GID>141</GID>
<name>N_in0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71,-29.5,74.5,-29.5</points>
<connection>
<GID>173</GID>
<name>OUT</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire></page 9></circuit>