<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>12.9741,-7.575,104.926,-53.025</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>29.5,-10.5</position>
<gparam>LABEL_TEXT Y=(A+B')(B+C')</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_INVERTER</type>
<position>34.5,-20.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>23,-18.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>22.5,-21</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AE_OR2</type>
<position>43.5,-20.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>38,-17</position>
<gparam>LABEL_TEXT B'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_TOGGLE</type>
<position>31,-29.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>30,-32</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AE_OR2</type>
<position>47,-40.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_INVERTER</type>
<position>34.5,-40.5</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_AND2</type>
<position>62.5,-20</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>24,-40.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>23.5,-43</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>41,-36.5</position>
<gparam>LABEL_TEXT C'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>38,-49</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>35,-48.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>GA_LED</type>
<position>63.5,-25.5</position>
<input>
<ID>N_in3</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>53.5,-16.5</position>
<gparam>LABEL_TEXT (A+B')</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>57.5,-42.5</position>
<gparam>LABEL_TEXT (B+C')</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_LABEL</type>
<position>63.5,-28</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-20.5,28,-18.5</points>
<intersection>-20.5 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-20.5,31.5,-20.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-18.5,28,-18.5</points>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-20.5,39,-19.5</points>
<intersection>-20.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-19.5,40.5,-19.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-20.5,39,-20.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-29.5,36.5,-21.5</points>
<intersection>-29.5 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-29.5,36.5,-29.5</points>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-21.5,40.5,-21.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-20.5,48,-19</points>
<intersection>-20.5 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-19,59.5,-19</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-20.5,48,-20.5</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-40.5,40.5,-39.5</points>
<intersection>-40.5 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-39.5,44,-39.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-40.5,40.5,-40.5</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-40.5,31.5,-40.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-49,42,-41.5</points>
<intersection>-49 2</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-41.5,44,-41.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>42 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-49,42,-49</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-40.5,58.5,-21</points>
<intersection>-40.5 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-21,59.5,-21</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>58.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>50,-40.5,58.5,-40.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>58.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-24.5,75,-20</points>
<intersection>-24.5 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-20,75,-20</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63.5,-24.5,75,-24.5</points>
<connection>
<GID>46</GID>
<name>N_in3</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-12.3472,24.1784,79.6046,-21.2716</PageViewport>
<gate>
<ID>3</ID>
<type>AE_OR3</type>
<position>41,11.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<input>
<ID>IN_2</ID>8 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>2,27</position>
<gparam>LABEL_TEXT F=AC+BC'+A'BC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_AND2</type>
<position>8.5,15</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_TOGGLE</type>
<position>-4,17.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>-3.5,12.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>-7,18</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>-7,13</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>7,11.5</position>
<gparam>LABEL_TEXT AC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_INVERTER</type>
<position>-2,3</position>
<input>
<ID>IN_0</ID>21 </input>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_TOGGLE</type>
<position>-10,5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>-10,2</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>AA_AND2</type>
<position>9,3</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>3,6</position>
<gparam>LABEL_TEXT C'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>-2,-5.5</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>-2,-2</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>8,-1.5</position>
<gparam>LABEL_TEXT BC'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_AND3</type>
<position>39.5,-13.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>26 </input>
<input>
<ID>IN_2</ID>25 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>20,-17</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_TOGGLE</type>
<position>20,-12.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_INVERTER</type>
<position>18,-7.5</position>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_TOGGLE</type>
<position>10,-7.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>25,-5</position>
<gparam>LABEL_TEXT A'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>17,-12</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>16.5,-16.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>GA_LED</type>
<position>60,8</position>
<input>
<ID>N_in3</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AA_LABEL</type>
<position>35.5,-6.5</position>
<gparam>LABEL_TEXT A'BC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_LABEL</type>
<position>45.5,17</position>
<gparam>LABEL_TEXT AC+BC'+A'BC</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>60,5.5</position>
<gparam>LABEL_TEXT F</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,9,60,11.5</points>
<connection>
<GID>112</GID>
<name>N_in3</name></connection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44,11.5,60,11.5</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,13.5,19.5,15</points>
<intersection>13.5 1</intersection>
<intersection>15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,13.5,38,13.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,15,19.5,15</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,3,19.5,11.5</points>
<intersection>3 2</intersection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,11.5,38,11.5</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,3,19.5,3</points>
<connection>
<GID>82</GID>
<name>OUT</name></connection>
<intersection>19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-13.5,37.5,9.5</points>
<intersection>-13.5 2</intersection>
<intersection>9.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-13.5,42.5,-13.5</points>
<connection>
<GID>92</GID>
<name>OUT</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>37.5,9.5,38,9.5</points>
<connection>
<GID>3</GID>
<name>IN_2</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1.5,16,1.5,17.5</points>
<intersection>16 1</intersection>
<intersection>17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1.5,16,5.5,16</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-2,17.5,1.5,17.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,12.5,2,14</points>
<intersection>12.5 2</intersection>
<intersection>14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,14,5.5,14</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-1.5,12.5,2,12.5</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6.5,3,-6.5,5</points>
<intersection>3 1</intersection>
<intersection>5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-6.5,3,-5,3</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>-6.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,5,-6.5,5</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>-6.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3.5,3,3.5,4</points>
<intersection>3 2</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3.5,4,6,4</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<intersection>3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1,3,3.5,3</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>3,-5.5,3,2</points>
<intersection>-5.5 2</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,2,6,2</points>
<connection>
<GID>82</GID>
<name>IN_1</name></connection>
<intersection>3 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>0,-5.5,3,-5.5</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>3 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-15.5,36.5,-15.5</points>
<connection>
<GID>92</GID>
<name>IN_2</name></connection>
<intersection>22 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22,-17,22,-15.5</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>-15.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>22,-13.5,36.5,-13.5</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<intersection>22 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22,-13.5,22,-12.5</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>-13.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,-7.5,15,-7.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-11.5,29,-7.5</points>
<intersection>-11.5 1</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-11.5,36.5,-11.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>21,-7.5,29,-7.5</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-0.101156,6.00992,122.501,-54.5901</PageViewport>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>56.5,-7</position>
<gparam>LABEL_TEXT DLD LAB PROJECT</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>56,-16</position>
<gparam>LABEL_TEXT TOPIC: REGISTER SHIFT: LEFT-RIGHT</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>56,-25</position>
<gparam>LABEL_TEXT NAME: ALI AKBER</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>55,-33.5</position>
<gparam>LABEL_TEXT ROLL NO: R036</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate></page 2>
<page 3>
<PageViewport>-0.101156,1.711e-006,122.501,-60.6</PageViewport></page 3>
<page 4>
<PageViewport>-0.101156,1.711e-006,122.501,-60.6</PageViewport></page 4>
<page 5>
<PageViewport>-0.101156,1.711e-006,122.501,-60.6</PageViewport></page 5>
<page 6>
<PageViewport>-0.101156,1.711e-006,122.501,-60.6</PageViewport></page 6>
<page 7>
<PageViewport>-0.101156,1.711e-006,122.501,-60.6</PageViewport></page 7>
<page 8>
<PageViewport>-0.101156,1.711e-006,122.501,-60.6</PageViewport></page 8>
<page 9>
<PageViewport>-0.101156,1.711e-006,122.501,-60.6</PageViewport></page 9></circuit>