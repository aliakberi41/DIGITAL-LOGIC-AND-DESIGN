<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-15,-6,107.4,-66.5</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>37.5,-11</position>
<gparam>LABEL_TEXT SHIFT RIGHT REGISTERS</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>77,-10.5</position>
<gparam>LABEL_TEXT (SISO)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AE_DFF_LOW_NT</type>
<position>-55,-14</position>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>21</ID>
<type>AE_DFF_LOW</type>
<position>20,-24</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT_0</ID>11 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>23</ID>
<type>AE_DFF_LOW</type>
<position>35,-24.5</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT_0</ID>12 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>25</ID>
<type>AE_DFF_LOW</type>
<position>49.5,-23</position>
<input>
<ID>IN_0</ID>12 </input>
<output>
<ID>OUT_0</ID>13 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>27</ID>
<type>AE_DFF_LOW</type>
<position>63.5,-24</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>14 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_TOGGLE</type>
<position>-0.5,-18.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>74.5,-22</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>BB_CLOCK</type>
<position>-1.5,-31.5</position>
<output>
<ID>CLK</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14,-39,14,-25</points>
<intersection>-39 1</intersection>
<intersection>-31.5 17</intersection>
<intersection>-25 7</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14,-39,60.5,-39</points>
<intersection>14 0</intersection>
<intersection>32 6</intersection>
<intersection>46.5 5</intersection>
<intersection>60.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>60.5,-39,60.5,-25</points>
<connection>
<GID>27</GID>
<name>clock</name></connection>
<intersection>-39 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>46.5,-39,46.5,-24</points>
<connection>
<GID>25</GID>
<name>clock</name></connection>
<intersection>-39 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>32,-39,32,-25.5</points>
<connection>
<GID>23</GID>
<name>clock</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>14,-25,17,-25</points>
<connection>
<GID>21</GID>
<name>clock</name></connection>
<intersection>14 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>2.5,-31.5,14,-31.5</points>
<connection>
<GID>50</GID>
<name>CLK</name></connection>
<intersection>14 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>9,-22,9,-18.5</points>
<intersection>-22 1</intersection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-22,17,-22</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>9 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1.5,-18.5,9,-18.5</points>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection>
<intersection>9 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-22.5,27.5,-22</points>
<intersection>-22.5 1</intersection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-22.5,32,-22.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-22,27.5,-22</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-22.5,42,-21</points>
<intersection>-22.5 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-21,46.5,-21</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>42 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-22.5,42,-22.5</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-22,56.5,-21</points>
<intersection>-22 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-22,60.5,-22</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52.5,-21,56.5,-21</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>66.5,-22,73.5,-22</points>
<connection>
<GID>48</GID>
<name>N_in0</name></connection>
<connection>
<GID>27</GID>
<name>OUT_0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-3,6,119.4,-54.5</PageViewport>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>48,2.5</position>
<gparam>LABEL_TEXT SHIFT LEFT REGISTER</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>84.5,2.5</position>
<gparam>LABEL_TEXT (SISO)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AE_DFF_LOW</type>
<position>82,-25.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>6 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_DFF_LOW</type>
<position>61.5,-25.5</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>7 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>12</ID>
<type>AE_DFF_LOW</type>
<position>41,-25.5</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>9 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_DFF_LOW</type>
<position>23.5,-25.5</position>
<input>
<ID>IN_0</ID>9 </input>
<output>
<ID>OUT_0</ID>15 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>95.5,-29</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>BB_CLOCK</type>
<position>92.5,-18.5</position>
<output>
<ID>CLK</ID>4 </output>
<gparam>angle 180</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>9,-23.5</position>
<input>
<ID>N_in1</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-13,88.5,-13</points>
<intersection>26.5 9</intersection>
<intersection>44 7</intersection>
<intersection>64.5 4</intersection>
<intersection>85 5</intersection>
<intersection>88.5 10</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>64.5,-24.5,64.5,-13</points>
<connection>
<GID>10</GID>
<name>clock</name></connection>
<intersection>-13 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>85,-24.5,85,-13</points>
<connection>
<GID>8</GID>
<name>clock</name></connection>
<intersection>-13 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>44,-24.5,44,-13</points>
<connection>
<GID>12</GID>
<name>clock</name></connection>
<intersection>-13 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>26.5,-24.5,26.5,-13</points>
<connection>
<GID>14</GID>
<name>clock</name></connection>
<intersection>-13 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>88.5,-18.5,88.5,-13</points>
<connection>
<GID>19</GID>
<name>CLK</name></connection>
<intersection>-13 1</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-29,89,-27.5</points>
<intersection>-29 2</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-27.5,89,-27.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89,-29,93.5,-29</points>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64.5,-27.5,79,-27.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>44,-27.5,58.5,-27.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-27.5,38,-27.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-27.5,15,-23.5</points>
<intersection>-27.5 2</intersection>
<intersection>-23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-23.5,15,-23.5</points>
<connection>
<GID>22</GID>
<name>N_in1</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,-27.5,20.5,-27.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-6,6,116.4,-54.5</PageViewport>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>46.5,2</position>
<gparam>LABEL_TEXT RIGHT SHIFT REGISTER</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>82.5,2</position>
<gparam>LABEL_TEXT (SIPO)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AE_DFF_LOW</type>
<position>22.5,-23</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>3 </output>
<input>
<ID>clock</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>16</ID>
<type>AE_DFF_LOW</type>
<position>39.5,-23</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>16 </output>
<input>
<ID>clock</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_DFF_LOW</type>
<position>57,-23</position>
<input>
<ID>IN_0</ID>16 </input>
<output>
<ID>OUT_0</ID>17 </output>
<input>
<ID>clock</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_DFF_LOW</type>
<position>80,-23</position>
<input>
<ID>IN_0</ID>17 </input>
<output>
<ID>OUT_0</ID>18 </output>
<input>
<ID>clock</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_TOGGLE</type>
<position>9.5,-16</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>31</ID>
<type>BB_CLOCK</type>
<position>6,-24</position>
<output>
<ID>CLK</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>33</ID>
<type>GA_LED</type>
<position>91,-23</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>GA_LED</type>
<position>28,-9</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>GA_LED</type>
<position>44.5,-9</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>GA_LED</type>
<position>62,-9</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-21,15.5,-16</points>
<intersection>-21 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,-21,19.5,-21</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-16,15.5,-16</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-33.5,77,-33.5</points>
<intersection>10 6</intersection>
<intersection>19.5 5</intersection>
<intersection>35 8</intersection>
<intersection>54 7</intersection>
<intersection>77 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>77,-33.5,77,-24</points>
<connection>
<GID>26</GID>
<name>clock</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>19.5,-33.5,19.5,-24</points>
<connection>
<GID>11</GID>
<name>clock</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>10,-33.5,10,-24</points>
<connection>
<GID>31</GID>
<name>CLK</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>54,-33.5,54,-24</points>
<connection>
<GID>20</GID>
<name>clock</name></connection>
<intersection>-33.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>35,-33.5,35,-24</points>
<intersection>-33.5 1</intersection>
<intersection>-24 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>35,-24,36.5,-24</points>
<connection>
<GID>16</GID>
<name>clock</name></connection>
<intersection>35 8</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25.5,-21,36.5,-21</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>30.5 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>30.5,-21,30.5,-9</points>
<intersection>-21 1</intersection>
<intersection>-9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>27,-9,30.5,-9</points>
<connection>
<GID>35</GID>
<name>N_in0</name></connection>
<intersection>30.5 2</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>42.5,-21,54,-21</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<connection>
<GID>16</GID>
<name>OUT_0</name></connection>
<intersection>47.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47.5,-21,47.5,-9</points>
<intersection>-21 1</intersection>
<intersection>-9 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>43.5,-9,47.5,-9</points>
<connection>
<GID>37</GID>
<name>N_in0</name></connection>
<intersection>47.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>60,-21,77,-21</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>64 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>64,-21,64,-9</points>
<intersection>-21 1</intersection>
<intersection>-9 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>61,-9,64,-9</points>
<connection>
<GID>39</GID>
<name>N_in0</name></connection>
<intersection>64 3</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-23,86.5,-21</points>
<intersection>-23 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-23,90,-23</points>
<connection>
<GID>33</GID>
<name>N_in0</name></connection>
<intersection>86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83,-21,86.5,-21</points>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,7.54211e-007,122.4,-60.5</PageViewport>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>55.5,-3.5</position>
<gparam>LABEL_TEXT LEFT SHIFT REGISTER</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>91,-3.5</position>
<gparam>LABEL_TEXT (SIPO)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AE_DFF_LOW</type>
<position>19,-26</position>
<input>
<ID>IN_0</ID>24 </input>
<output>
<ID>OUT_0</ID>25 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>49</ID>
<type>AE_DFF_LOW</type>
<position>36,-25.5</position>
<input>
<ID>IN_0</ID>23 </input>
<output>
<ID>OUT_0</ID>24 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>52</ID>
<type>AE_DFF_LOW</type>
<position>55.5,-25.5</position>
<input>
<ID>IN_0</ID>22 </input>
<output>
<ID>OUT_0</ID>23 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>54</ID>
<type>AE_DFF_LOW</type>
<position>71,-25</position>
<input>
<ID>IN_0</ID>21 </input>
<output>
<ID>OUT_0</ID>22 </output>
<input>
<ID>clock</ID>20 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>88,-31.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>60</ID>
<type>BB_CLOCK</type>
<position>87,-20.5</position>
<output>
<ID>CLK</ID>20 </output>
<gparam>angle 180</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>8,-26.5</position>
<input>
<ID>N_in1</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>GA_LED</type>
<position>32.5,-41</position>
<input>
<ID>N_in3</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>GA_LED</type>
<position>52.5,-41.5</position>
<input>
<ID>N_in3</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>GA_LED</type>
<position>68,-42</position>
<input>
<ID>N_in3</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-20.5,78.5,-14</points>
<intersection>-20.5 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-14,78.5,-14</points>
<intersection>22 9</intersection>
<intersection>39 7</intersection>
<intersection>58.5 5</intersection>
<intersection>74 3</intersection>
<intersection>78.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78.5,-20.5,83,-20.5</points>
<connection>
<GID>60</GID>
<name>CLK</name></connection>
<intersection>78.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74,-24,74,-14</points>
<connection>
<GID>54</GID>
<name>clock</name></connection>
<intersection>-14 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>58.5,-24.5,58.5,-14</points>
<connection>
<GID>52</GID>
<name>clock</name></connection>
<intersection>-14 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>39,-24.5,39,-14</points>
<connection>
<GID>49</GID>
<name>clock</name></connection>
<intersection>-14 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>22,-25,22,-14</points>
<connection>
<GID>45</GID>
<name>clock</name></connection>
<intersection>-14 1</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-31.5,80,-27</points>
<intersection>-31.5 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-27,80,-27</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80,-31.5,86,-31.5</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-27.5,63,-27</points>
<intersection>-27.5 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>58.5,-27.5,63,-27.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>63,-27,68,-27</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>63 0</intersection>
<intersection>68 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>68,-41,68,-27</points>
<connection>
<GID>68</GID>
<name>N_in3</name></connection>
<intersection>-27 2</intersection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-27.5,52.5,-27.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>52.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>52.5,-40.5,52.5,-27.5</points>
<connection>
<GID>66</GID>
<name>N_in3</name></connection>
<intersection>-27.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-28,27.5,-27.5</points>
<intersection>-28 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-28,27.5,-28</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-27.5,33,-27.5</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>27.5 0</intersection>
<intersection>32.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32.5,-40,32.5,-27.5</points>
<connection>
<GID>64</GID>
<name>N_in3</name></connection>
<intersection>-27.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-28,12.5,-26.5</points>
<intersection>-28 2</intersection>
<intersection>-26.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-26.5,12.5,-26.5</points>
<connection>
<GID>62</GID>
<name>N_in1</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-28,16,-28</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>-12,7.54211e-007,110.4,-60.5</PageViewport>
<gate>
<ID>9</ID>
<type>AE_DFF_LOW</type>
<position>29,-46</position>
<input>
<ID>IN_0</ID>26 </input>
<output>
<ID>OUT_0</ID>30 </output>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>18</ID>
<type>AE_DFF_LOW</type>
<position>46,-46</position>
<input>
<ID>IN_0</ID>33 </input>
<output>
<ID>OUT_0</ID>35 </output>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>28</ID>
<type>AE_DFF_LOW</type>
<position>66,-46</position>
<input>
<ID>IN_0</ID>38 </input>
<output>
<ID>OUT_0</ID>40 </output>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>32</ID>
<type>AE_DFF_LOW</type>
<position>85,-45.5</position>
<input>
<ID>IN_0</ID>43 </input>
<output>
<ID>OUT_0</ID>44 </output>
<input>
<ID>clock</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>22.5,-8.5</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>41.5,-9</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>60.5,-7</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>80.5,-8.5</position>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>55</ID>
<type>BB_CLOCK</type>
<position>11,-51.5</position>
<output>
<ID>CLK</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_AND2</type>
<position>29.5,-18.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_AND2</type>
<position>36,-18.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_AND2</type>
<position>49,-17.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_AND2</type>
<position>56,-17.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>41,-2</position>
<gparam>LABEL_TEXT RIGHT SHIFT REGISTER </gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>77,-2</position>
<gparam>LABEL_TEXT (PISO)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_AND2</type>
<position>70,-20</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_AND2</type>
<position>76.5,-19.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_INVERTER</type>
<position>6,-15</position>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_TOGGLE</type>
<position>-2.5,-14.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>83</ID>
<type>AE_OR2</type>
<position>34,-27.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>AE_OR2</type>
<position>53,-26.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>87</ID>
<type>AE_OR2</type>
<position>74,-28</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>89</ID>
<type>GA_LED</type>
<position>96.5,-43.5</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-54,20.5,-51.5</points>
<intersection>-54 1</intersection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-54,82,-54</points>
<intersection>20.5 0</intersection>
<intersection>26 5</intersection>
<intersection>43 4</intersection>
<intersection>63 7</intersection>
<intersection>82 9</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>15,-51.5,20.5,-51.5</points>
<connection>
<GID>55</GID>
<name>CLK</name></connection>
<intersection>20.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>43,-54,43,-47</points>
<connection>
<GID>18</GID>
<name>clock</name></connection>
<intersection>-54 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>26,-54,26,-47</points>
<connection>
<GID>9</GID>
<name>clock</name></connection>
<intersection>-54 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>63,-54,63,-47</points>
<connection>
<GID>28</GID>
<name>clock</name></connection>
<intersection>-54 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>82,-54,82,-46.5</points>
<connection>
<GID>32</GID>
<name>clock</name></connection>
<intersection>-54 1</intersection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-44,22.5,-10.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-44,26,-44</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-11.5,71,-11.5</points>
<intersection>-0.5 3</intersection>
<intersection>3 5</intersection>
<intersection>30.5 4</intersection>
<intersection>50 7</intersection>
<intersection>71 9</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-0.5,-14.5,-0.5,-11.5</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>30.5,-15.5,30.5,-11.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>3,-15,3,-11.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>50,-14.5,50,-11.5</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>71,-17,71,-11.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>-11.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-15.5,37,-14</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>-14 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>41.5,-14,41.5,-11</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>37,-14,41.5,-14</points>
<intersection>37 0</intersection>
<intersection>41.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-15.5,35,-13</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>9,-13,75.5,-13</points>
<intersection>9 2</intersection>
<intersection>35 0</intersection>
<intersection>55 4</intersection>
<intersection>75.5 6</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>9,-15,9,-13</points>
<connection>
<GID>79</GID>
<name>OUT_0</name></connection>
<intersection>-13 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>55,-14.5,55,-13</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>-13 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>75.5,-16.5,75.5,-13</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>-13 1</intersection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-40,25.5,-15.5</points>
<intersection>-40 1</intersection>
<intersection>-15.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-40,32,-40</points>
<intersection>25.5 0</intersection>
<intersection>32 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>32,-44,32,-40</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>25.5,-15.5,28.5,-15.5</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-24.5,33,-21.5</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-21.5,33,-21.5</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-24.5,35,-23</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>-23 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>40,-23,40,-21.5</points>
<intersection>-23 2</intersection>
<intersection>-21.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35,-23,40,-23</points>
<intersection>35 0</intersection>
<intersection>40 1</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>36,-21.5,40,-21.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>40 1</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-44,34,-30.5</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-44,43,-44</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-14.5,60.5,-9</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>57,-14.5,60.5,-14.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-41,43,-14.5</points>
<intersection>-41 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-41,49,-41</points>
<intersection>43 0</intersection>
<intersection>49 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>43,-14.5,48,-14.5</points>
<connection>
<GID>65</GID>
<name>IN_1</name></connection>
<intersection>43 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49,-44,49,-41</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>-41 1</intersection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-23.5,52,-22</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>-22 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>49,-22,49,-20.5</points>
<connection>
<GID>65</GID>
<name>OUT</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>49,-22,52,-22</points>
<intersection>49 1</intersection>
<intersection>52 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-23.5,54,-22</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>-22 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>56,-22,56,-20.5</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>54,-22,56,-22</points>
<intersection>54 0</intersection>
<intersection>56 1</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53,-44,53,-29.5</points>
<connection>
<GID>85</GID>
<name>OUT</name></connection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-44,63,-44</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>53 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-16.5,77.5,-12</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>-12 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>80.5,-12,80.5,-10.5</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-12,80.5,-12</points>
<intersection>77.5 0</intersection>
<intersection>80.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-41,64.5,-17</points>
<intersection>-41 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64.5,-17,69,-17</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-41,69,-41</points>
<intersection>64.5 0</intersection>
<intersection>69 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>69,-44,69,-41</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>-41 2</intersection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-25,73,-24</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<intersection>-24 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>70,-24,70,-23</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>70,-24,73,-24</points>
<intersection>70 1</intersection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-25,75,-23.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>-23.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>76.5,-23.5,76.5,-22.5</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>75,-23.5,76.5,-23.5</points>
<intersection>75 0</intersection>
<intersection>76.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74,-43.5,74,-31</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,-43.5,82,-43.5</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>74 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-43.5,95.5,-43.5</points>
<connection>
<GID>89</GID>
<name>N_in0</name></connection>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>0,3,122.4,-57.5</PageViewport>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>52,1</position>
<gparam>LABEL_TEXT LEFT SHIFT REGISTER</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>85,1</position>
<gparam>LABEL_TEXT (PISO)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AE_DFF_LOW</type>
<position>89,-44.5</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUTINV_0</ID>50 </output>
<input>
<ID>clock</ID>46 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>93</ID>
<type>AE_DFF_LOW</type>
<position>66.5,-44.5</position>
<input>
<ID>IN_0</ID>55 </input>
<output>
<ID>OUTINV_0</ID>56 </output>
<input>
<ID>clock</ID>46 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>95</ID>
<type>AE_DFF_LOW</type>
<position>44.5,-44.5</position>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUTINV_0</ID>66 </output>
<input>
<ID>clock</ID>46 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>97</ID>
<type>AE_DFF_LOW</type>
<position>24.5,-44.5</position>
<input>
<ID>IN_0</ID>63 </input>
<output>
<ID>OUTINV_0</ID>67 </output>
<input>
<ID>clock</ID>46 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>99</ID>
<type>GA_LED</type>
<position>6.5,-43</position>
<input>
<ID>N_in1</ID>67 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>BB_CLOCK</type>
<position>103.5,-45.5</position>
<output>
<ID>CLK</ID>46 </output>
<gparam>angle 180</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_TOGGLE</type>
<position>30.5,-6</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_TOGGLE</type>
<position>52.5,-4</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_TOGGLE</type>
<position>73.5,-4.5</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_TOGGLE</type>
<position>112,-11</position>
<output>
<ID>OUT_0</ID>47 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_INVERTER</type>
<position>101.5,-11.5</position>
<input>
<ID>IN_0</ID>47 </input>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_AND2</type>
<position>33,-17.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>65 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AA_AND2</type>
<position>39,-17.5</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AE_OR2</type>
<position>36.5,-25</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>AA_AND2</type>
<position>53,-18</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_AND2</type>
<position>59.5,-18</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>AE_OR2</type>
<position>56.5,-26</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_AND2</type>
<position>75.5,-18</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_AND2</type>
<position>82,-18</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>131</ID>
<type>AE_OR2</type>
<position>79.5,-26</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_TOGGLE</type>
<position>92.5,-4.5</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-54,95.5,-45.5</points>
<intersection>-54 1</intersection>
<intersection>-45.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-54,95.5,-54</points>
<intersection>29 9</intersection>
<intersection>49.5 7</intersection>
<intersection>71.5 4</intersection>
<intersection>93.5 5</intersection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,-45.5,99.5,-45.5</points>
<connection>
<GID>101</GID>
<name>CLK</name></connection>
<intersection>95.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>71.5,-54,71.5,-43.5</points>
<intersection>-54 1</intersection>
<intersection>-43.5 11</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>93.5,-54,93.5,-43.5</points>
<intersection>-54 1</intersection>
<intersection>-43.5 10</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>49.5,-54,49.5,-43.5</points>
<intersection>-54 1</intersection>
<intersection>-43.5 12</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>29,-54,29,-43.5</points>
<intersection>-54 1</intersection>
<intersection>-43.5 13</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>92,-43.5,93.5,-43.5</points>
<connection>
<GID>91</GID>
<name>clock</name></connection>
<intersection>93.5 5</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>69.5,-43.5,71.5,-43.5</points>
<connection>
<GID>93</GID>
<name>clock</name></connection>
<intersection>71.5 4</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>47.5,-43.5,49.5,-43.5</points>
<connection>
<GID>95</GID>
<name>clock</name></connection>
<intersection>49.5 7</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>27.5,-43.5,29,-43.5</points>
<connection>
<GID>97</GID>
<name>clock</name></connection>
<intersection>29 9</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-11,107,-8</points>
<intersection>-11 2</intersection>
<intersection>-8 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38,-8,107,-8</points>
<intersection>38 8</intersection>
<intersection>58.5 6</intersection>
<intersection>81 3</intersection>
<intersection>104.5 4</intersection>
<intersection>107 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>107,-11,110,-11</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<intersection>107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>81,-15,81,-8</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>-8 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>104.5,-11.5,104.5,-8</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-8 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>58.5,-15,58.5,-8</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>-8 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>38,-14.5,38,-8</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>-8 1</intersection></vsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-46.5,92.5,-6.5</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,-46.5,92.5,-46.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-43.5,85.5,-15</points>
<intersection>-43.5 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-43.5,86,-43.5</points>
<connection>
<GID>91</GID>
<name>OUTINV_0</name></connection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>83,-15,85.5,-15</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-15,76.5,-10.5</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-10.5,98.5,-10.5</points>
<intersection>34 6</intersection>
<intersection>54 3</intersection>
<intersection>76.5 0</intersection>
<intersection>98.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54,-15,54,-10.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>98.5,-11.5,98.5,-10.5</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<intersection>-10.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>34,-14.5,34,-10.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>-10.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-15,74.5,-12</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<intersection>-12 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>73.5,-12,73.5,-6.5</points>
<connection>
<GID>107</GID>
<name>OUT_0</name></connection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-12,74.5,-12</points>
<intersection>73.5 1</intersection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-23,78.5,-22</points>
<connection>
<GID>131</GID>
<name>IN_1</name></connection>
<intersection>-22 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>75.5,-22,75.5,-21</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>75.5,-22,78.5,-22</points>
<intersection>75.5 1</intersection>
<intersection>78.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-23,80.5,-22</points>
<connection>
<GID>131</GID>
<name>IN_0</name></connection>
<intersection>-22 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>82,-22,82,-21</points>
<connection>
<GID>129</GID>
<name>OUT</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>80.5,-22,82,-22</points>
<intersection>80.5 0</intersection>
<intersection>82 1</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-46.5,79.5,-29</points>
<connection>
<GID>131</GID>
<name>OUT</name></connection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-46.5,79.5,-46.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63,-43.5,63,-15</points>
<intersection>-43.5 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63,-43.5,63.5,-43.5</points>
<connection>
<GID>93</GID>
<name>OUTINV_0</name></connection>
<intersection>63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60.5,-15,63,-15</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>63 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-15,52,-11.5</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>52.5,-11.5,52.5,-6</points>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>52,-11.5,52.5,-11.5</points>
<intersection>52 0</intersection>
<intersection>52.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-23,55.5,-22</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>-22 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>53,-22,53,-21</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>53,-22,55.5,-22</points>
<intersection>53 1</intersection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>57.5,-23,57.5,-22</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>-22 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>59.5,-22,59.5,-21</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57.5,-22,59.5,-22</points>
<intersection>57.5 0</intersection>
<intersection>59.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-46.5,56.5,-29</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47.5,-46.5,56.5,-46.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-22,35.5,-21</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>-21 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>33,-21,33,-20.5</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>33,-21,35.5,-21</points>
<intersection>33 1</intersection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-22,37.5,-21</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>-21 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>39,-21,39,-20.5</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>37.5,-21,39,-21</points>
<intersection>37.5 0</intersection>
<intersection>39 1</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-46.5,36.5,-28</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-46.5,36.5,-46.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>36.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-14.5,32,-11</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>-11 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>30.5,-11,30.5,-8</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>-11 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-11,32,-11</points>
<intersection>30.5 1</intersection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-43.5,41.5,-14.5</points>
<connection>
<GID>95</GID>
<name>OUTINV_0</name></connection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>40,-14.5,41.5,-14.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-43.5,14.5,-43</points>
<intersection>-43.5 1</intersection>
<intersection>-43 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-43.5,21.5,-43.5</points>
<connection>
<GID>97</GID>
<name>OUTINV_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-43,14.5,-43</points>
<connection>
<GID>99</GID>
<name>N_in1</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>0,7.54211e-007,122.4,-60.5</PageViewport>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>57,-3</position>
<gparam>LABEL_TEXT SHIFT RIGHT REGISTER</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>92.5,-3</position>
<gparam>LABEL_TEXT (PIPO)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AE_DFF_LOW</type>
<position>25,-30</position>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>48 </output>
<input>
<ID>clock</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>63</ID>
<type>AE_DFF_LOW</type>
<position>42,-29.5</position>
<input>
<ID>IN_0</ID>72 </input>
<output>
<ID>OUT_0</ID>64 </output>
<input>
<ID>clock</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>71</ID>
<type>AE_DFF_LOW</type>
<position>59.5,-30</position>
<input>
<ID>IN_0</ID>73 </input>
<output>
<ID>OUT_0</ID>68 </output>
<input>
<ID>clock</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>78</ID>
<type>AE_DFF_LOW</type>
<position>76,-29</position>
<input>
<ID>IN_0</ID>74 </input>
<output>
<ID>OUT_0</ID>70 </output>
<input>
<ID>clock</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>82</ID>
<type>GA_LED</type>
<position>31.5,-46</position>
<input>
<ID>N_in3</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>GA_LED</type>
<position>49.5,-46</position>
<input>
<ID>N_in3</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>GA_LED</type>
<position>66,-46</position>
<input>
<ID>N_in3</ID>68 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_TOGGLE</type>
<position>24,-10</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_TOGGLE</type>
<position>41.5,-10</position>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_TOGGLE</type>
<position>59,-9.5</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_TOGGLE</type>
<position>76,-9.5</position>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>112</ID>
<type>BB_CLOCK</type>
<position>8,-35</position>
<output>
<ID>CLK</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>116</ID>
<type>GA_LED</type>
<position>87,-47</position>
<input>
<ID>N_in3</ID>70 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17,-37.5,17,-35</points>
<intersection>-37.5 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,-37.5,73,-37.5</points>
<intersection>17 0</intersection>
<intersection>22 4</intersection>
<intersection>39 3</intersection>
<intersection>56.5 6</intersection>
<intersection>73 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-35,17,-35</points>
<connection>
<GID>112</GID>
<name>CLK</name></connection>
<intersection>17 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>39,-37.5,39,-30.5</points>
<connection>
<GID>63</GID>
<name>clock</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>22,-37.5,22,-31</points>
<connection>
<GID>57</GID>
<name>clock</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>56.5,-37.5,56.5,-31</points>
<connection>
<GID>71</GID>
<name>clock</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>73,-37.5,73,-30</points>
<connection>
<GID>78</GID>
<name>clock</name></connection>
<intersection>-37.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-45,31.5,-28</points>
<connection>
<GID>82</GID>
<name>N_in3</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-28,31.5,-28</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-45,49.5,-27.5</points>
<connection>
<GID>86</GID>
<name>N_in3</name></connection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-27.5,49.5,-27.5</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-45,66,-28</points>
<connection>
<GID>90</GID>
<name>N_in3</name></connection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-28,66,-28</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>66 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-46,87,-27</points>
<connection>
<GID>116</GID>
<name>N_in3</name></connection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79,-27,87,-27</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-28,19.5,-16</points>
<intersection>-28 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>19.5,-28,22,-28</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-16,24,-16</points>
<intersection>19.5 0</intersection>
<intersection>24 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>24,-16,24,-12</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<intersection>-16 2</intersection></vsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-27.5,36.5,-16</points>
<intersection>-27.5 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36.5,-27.5,39,-27.5</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-16,41.5,-16</points>
<intersection>36.5 0</intersection>
<intersection>41.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>41.5,-16,41.5,-12</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<intersection>-16 2</intersection></vsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-28,54,-14.5</points>
<intersection>-28 1</intersection>
<intersection>-14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-28,56.5,-28</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-14.5,59,-14.5</points>
<intersection>54 0</intersection>
<intersection>59 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>59,-14.5,59,-11.5</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<intersection>-14.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-27,71.5,-11.5</points>
<intersection>-27 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-27,73,-27</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>71.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>71.5,-11.5,76,-11.5</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<intersection>71.5 0</intersection></hsegment></shape></wire></page 6>
<page 7>
<PageViewport>0,7.54211e-007,122.4,-60.5</PageViewport>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>56.5,-3</position>
<gparam>LABEL_TEXT SHIFT LEFT REGISTER</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>91.5,-3</position>
<gparam>LABEL_TEXT (PIPO)</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AE_DFF_LOW</type>
<position>22.5,-30.5</position>
<input>
<ID>IN_0</ID>76 </input>
<output>
<ID>OUT_0</ID>78 </output>
<input>
<ID>clock</ID>75 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>124</ID>
<type>AE_DFF_LOW</type>
<position>40,-30.5</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>84 </output>
<input>
<ID>clock</ID>75 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>128</ID>
<type>AE_DFF_LOW</type>
<position>56.5,-30</position>
<input>
<ID>IN_0</ID>85 </input>
<output>
<ID>OUT_0</ID>86 </output>
<input>
<ID>clock</ID>75 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>132</ID>
<type>AE_DFF_LOW</type>
<position>74.5,-30</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>88 </output>
<input>
<ID>clock</ID>75 </input>
<gparam>angle 180</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>135</ID>
<type>BB_CLOCK</type>
<position>90.5,-33</position>
<output>
<ID>CLK</ID>75 </output>
<gparam>angle 180</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>137</ID>
<type>AA_TOGGLE</type>
<position>26.5,-49.5</position>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>139</ID>
<type>GA_LED</type>
<position>16.5,-13.5</position>
<input>
<ID>N_in2</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>AA_TOGGLE</type>
<position>45,-51</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_TOGGLE</type>
<position>60.5,-50.5</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_TOGGLE</type>
<position>74,-52</position>
<output>
<ID>OUT_0</ID>87 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>147</ID>
<type>GA_LED</type>
<position>34,-12.5</position>
<input>
<ID>N_in2</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>GA_LED</type>
<position>50.5,-12.5</position>
<input>
<ID>N_in2</ID>86 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>151</ID>
<type>GA_LED</type>
<position>68,-11</position>
<input>
<ID>N_in2</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-42,82,-33</points>
<intersection>-42 1</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-42,82,-42</points>
<intersection>29 11</intersection>
<intersection>47.5 8</intersection>
<intersection>63 9</intersection>
<intersection>79 5</intersection>
<intersection>82 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-33,86.5,-33</points>
<connection>
<GID>135</GID>
<name>CLK</name></connection>
<intersection>82 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>79,-42,79,-29</points>
<intersection>-42 1</intersection>
<intersection>-29 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>77.5,-29,79,-29</points>
<connection>
<GID>132</GID>
<name>clock</name></connection>
<intersection>79 5</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>47.5,-42,47.5,-29.5</points>
<intersection>-42 1</intersection>
<intersection>-29.5 12</intersection></vsegment>
<vsegment>
<ID>9</ID>
<points>63,-42,63,-29</points>
<intersection>-42 1</intersection>
<intersection>-29 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>29,-42,29,-29.5</points>
<intersection>-42 1</intersection>
<intersection>-29.5 13</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>43,-29.5,47.5,-29.5</points>
<connection>
<GID>124</GID>
<name>clock</name></connection>
<intersection>47.5 8</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>25.5,-29.5,29,-29.5</points>
<connection>
<GID>120</GID>
<name>clock</name></connection>
<intersection>29 11</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>59.5,-29,63,-29</points>
<connection>
<GID>128</GID>
<name>clock</name></connection>
<intersection>63 9</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-47.5,26.5,-32.5</points>
<connection>
<GID>137</GID>
<name>OUT_0</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-32.5,26.5,-32.5</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>16.5,-32.5,16.5,-14.5</points>
<connection>
<GID>139</GID>
<name>N_in2</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16.5,-32.5,19.5,-32.5</points>
<connection>
<GID>120</GID>
<name>OUT_0</name></connection>
<intersection>16.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-49,45,-32.5</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43,-32.5,45,-32.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-32.5,34,-13.5</points>
<connection>
<GID>147</GID>
<name>N_in2</name></connection>
<intersection>-32.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-32.5,37,-32.5</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-48.5,60.5,-32</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59.5,-32,60.5,-32</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-32,50.5,-13.5</points>
<connection>
<GID>149</GID>
<name>N_in2</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-32,53.5,-32</points>
<connection>
<GID>128</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-49.5,77.5,-32</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>-49.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>74,-49.5,77.5,-49.5</points>
<intersection>74 3</intersection>
<intersection>77.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74,-50,74,-49.5</points>
<connection>
<GID>145</GID>
<name>OUT_0</name></connection>
<intersection>-49.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-32,68,-12</points>
<connection>
<GID>151</GID>
<name>N_in2</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-32,71.5,-32</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire></page 7>
<page 8>
<PageViewport>-3,3,119.4,-57.5</PageViewport>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>57.5,0</position>
<gparam>LABEL_TEXT BIDIRECTIONAL SHIFT REGISTER</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>5,-42</position>
<input>
<ID>N_in1</ID>100 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AE_DFF_LOW</type>
<position>23,-42.5</position>
<input>
<ID>IN_0</ID>82 </input>
<output>
<ID>OUT_0</ID>96 </output>
<input>
<ID>clear</ID>107 </input>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>59</ID>
<type>AE_DFF_LOW</type>
<position>46.5,-42</position>
<input>
<ID>IN_0</ID>100 </input>
<output>
<ID>OUT_0</ID>102 </output>
<input>
<ID>clear</ID>107 </input>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>75</ID>
<type>AE_DFF_LOW</type>
<position>72,-41</position>
<input>
<ID>IN_0</ID>101 </input>
<output>
<ID>OUT_0</ID>103 </output>
<input>
<ID>clear</ID>107 </input>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>84</ID>
<type>AE_DFF_LOW</type>
<position>99.5,-40.5</position>
<input>
<ID>IN_0</ID>99 </input>
<output>
<ID>OUT_0</ID>104 </output>
<input>
<ID>clear</ID>107 </input>
<input>
<ID>clock</ID>77 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>92</ID>
<type>AA_TOGGLE</type>
<position>1.5,-9</position>
<output>
<ID>OUT_0</ID>108 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_AND2</type>
<position>8,-19</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_AND2</type>
<position>15,-19</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>AE_OR2</type>
<position>12,-26.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_AND2</type>
<position>32,-18.5</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>90 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_AND2</type>
<position>40,-18</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>AE_OR2</type>
<position>36,-26</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>AA_AND2</type>
<position>57,-18</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_AND2</type>
<position>64.5,-18</position>
<input>
<ID>IN_0</ID>104 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>93 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>AE_OR2</type>
<position>61,-25.5</position>
<input>
<ID>IN_0</ID>93 </input>
<input>
<ID>IN_1</ID>92 </input>
<output>
<ID>OUT</ID>101 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_AND2</type>
<position>82.5,-17.5</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>94 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_AND2</type>
<position>89.5,-17.5</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>155</ID>
<type>AE_OR2</type>
<position>86,-25</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_INVERTER</type>
<position>13,-10.5</position>
<input>
<ID>IN_0</ID>108 </input>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>159</ID>
<type>BB_CLOCK</type>
<position>5.5,-49</position>
<output>
<ID>CLK</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_TOGGLE</type>
<position>0.5,-16</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>165</ID>
<type>AA_TOGGLE</type>
<position>96,-10</position>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 180</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>167</ID>
<type>GA_LED</type>
<position>106,-37.5</position>
<input>
<ID>N_in0</ID>104 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>AA_TOGGLE</type>
<position>5,-55</position>
<output>
<ID>OUT_0</ID>107 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>77</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>9.5,-49,96.5,-49</points>
<connection>
<GID>159</GID>
<name>CLK</name></connection>
<intersection>18 4</intersection>
<intersection>40 3</intersection>
<intersection>66 6</intersection>
<intersection>96.5 8</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>40,-49,40,-43</points>
<intersection>-49 1</intersection>
<intersection>-43 14</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>18,-49,18,-43.5</points>
<intersection>-49 1</intersection>
<intersection>-43.5 13</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>66,-49,66,-42</points>
<intersection>-49 1</intersection>
<intersection>-42 15</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>96.5,-49,96.5,-41.5</points>
<connection>
<GID>84</GID>
<name>clock</name></connection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>18,-43.5,20,-43.5</points>
<connection>
<GID>42</GID>
<name>clock</name></connection>
<intersection>18 4</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>40,-43,43.5,-43</points>
<connection>
<GID>59</GID>
<name>clock</name></connection>
<intersection>40 3</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>66,-42,69,-42</points>
<connection>
<GID>75</GID>
<name>clock</name></connection>
<intersection>66 6</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-23.5,11,-22.5</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>-22.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>8,-22.5,8,-22</points>
<connection>
<GID>96</GID>
<name>OUT</name></connection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>8,-22.5,11,-22.5</points>
<intersection>8 1</intersection>
<intersection>11 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-23.5,13,-22.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>-22.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>15,-22.5,15,-22</points>
<connection>
<GID>104</GID>
<name>OUT</name></connection>
<intersection>-22.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>13,-22.5,15,-22.5</points>
<intersection>13 0</intersection>
<intersection>15 1</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>3,-13.5,9,-13.5</points>
<intersection>3 3</intersection>
<intersection>9 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>9,-16,9,-13.5</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>-13.5 1</intersection></vsegment>
<vsegment>
<ID>3</ID>
<points>3,-16,3,-13.5</points>
<intersection>-16 4</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>2.5,-16,3,-16</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>3 3</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-40.5,12,-29.5</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<intersection>-40.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12,-40.5,20,-40.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>12 0</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-13.5,18.5,-7.5</points>
<intersection>-13.5 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>16,-7.5,88.5,-7.5</points>
<intersection>16 4</intersection>
<intersection>18.5 0</intersection>
<intersection>39 6</intersection>
<intersection>63.5 8</intersection>
<intersection>88.5 10</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>14,-13.5,18.5,-13.5</points>
<intersection>14 3</intersection>
<intersection>18.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14,-16,14,-13.5</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<intersection>-13.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>16,-10.5,16,-7.5</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>39,-15,39,-7.5</points>
<connection>
<GID>126</GID>
<name>IN_1</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>63.5,-15,63.5,-7.5</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>-7.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>88.5,-14.5,88.5,-7.5</points>
<connection>
<GID>153</GID>
<name>IN_1</name></connection>
<intersection>-7.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-23,35,-22</points>
<connection>
<GID>134</GID>
<name>IN_1</name></connection>
<intersection>-22 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>32,-22,32,-21.5</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>32,-22,35,-22</points>
<intersection>32 1</intersection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-23,37,-22</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>-22 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>40,-22,40,-21</points>
<connection>
<GID>126</GID>
<name>OUT</name></connection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>37,-22,40,-22</points>
<intersection>37 0</intersection>
<intersection>40 1</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-22.5,60,-21.5</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>57,-21.5,57,-21</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>57,-21.5,60,-21.5</points>
<intersection>57 1</intersection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62,-22.5,62,-21.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>64.5,-21.5,64.5,-21</points>
<connection>
<GID>142</GID>
<name>OUT</name></connection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>62,-21.5,64.5,-21.5</points>
<intersection>62 0</intersection>
<intersection>64.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-22,85,-21</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>-21 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>82.5,-21,82.5,-20.5</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-21,85,-21</points>
<intersection>82.5 1</intersection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-22,87,-21</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>-21 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>89.5,-21,89.5,-20.5</points>
<connection>
<GID>153</GID>
<name>OUT</name></connection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>87,-21,89.5,-21</points>
<intersection>87 0</intersection>
<intersection>89.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-42,27.5,-14</points>
<intersection>-42 1</intersection>
<intersection>-14 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-42,27.5,-42</points>
<intersection>26 5</intersection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-14,33,-14</points>
<intersection>27.5 0</intersection>
<intersection>33 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33,-15.5,33,-14</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>-14 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>26,-42,26,-40.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>-42 1</intersection></vsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-38.5,86,-28</points>
<connection>
<GID>155</GID>
<name>OUT</name></connection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,-38.5,96.5,-38.5</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-40,36,-29</points>
<connection>
<GID>134</GID>
<name>OUT</name></connection>
<intersection>-40 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>36,-40,43.5,-40</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>36 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-36,36,-36</points>
<intersection>5 3</intersection>
<intersection>36 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>5,-42,5,-36</points>
<intersection>-42 4</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>5,-42,6,-42</points>
<connection>
<GID>34</GID>
<name>N_in1</name></connection>
<intersection>5 3</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-39,61,-28.5</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-39,69,-39</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52,-40,52,-12.5</points>
<intersection>-40 1</intersection>
<intersection>-30.5 4</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-40,52,-40</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>52 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-12.5,58,-12.5</points>
<intersection>52 0</intersection>
<intersection>58 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>58,-15,58,-12.5</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20.5,-30.5,52,-30.5</points>
<intersection>20.5 5</intersection>
<intersection>52 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>20.5,-30.5,20.5,-16</points>
<intersection>-30.5 4</intersection>
<intersection>-16 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>16,-16,20.5,-16</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>20.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77,-39,77,-10.5</points>
<intersection>-39 1</intersection>
<intersection>-13 2</intersection>
<intersection>-10.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-39,77,-39</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>77 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-13,83.5,-13</points>
<intersection>77 0</intersection>
<intersection>83.5 5</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>41,-10.5,77,-10.5</points>
<intersection>41 4</intersection>
<intersection>77 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>41,-15,41,-10.5</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<intersection>-10.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>83.5,-14.5,83.5,-13</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>-13 2</intersection></vsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-34.5,71,-15</points>
<intersection>-34.5 1</intersection>
<intersection>-15 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-34.5,103,-34.5</points>
<intersection>71 0</intersection>
<intersection>103 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>103,-38.5,103,-34.5</points>
<intersection>-38.5 4</intersection>
<intersection>-37.5 5</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>65.5,-15,71,-15</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>102.5,-38.5,103,-38.5</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>103 2</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>103,-37.5,105,-37.5</points>
<connection>
<GID>167</GID>
<name>N_in0</name></connection>
<intersection>103 2</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-14.5,90.5,-10</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90.5,-10,94,-10</points>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-55,23,-46.5</points>
<connection>
<GID>42</GID>
<name>clear</name></connection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>7,-55,99.5,-55</points>
<connection>
<GID>171</GID>
<name>OUT_0</name></connection>
<intersection>23 0</intersection>
<intersection>46.5 3</intersection>
<intersection>72 5</intersection>
<intersection>99.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>46.5,-55,46.5,-46</points>
<connection>
<GID>59</GID>
<name>clear</name></connection>
<intersection>-55 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>72,-55,72,-45</points>
<connection>
<GID>75</GID>
<name>clear</name></connection>
<intersection>-55 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>99.5,-55,99.5,-44.5</points>
<connection>
<GID>84</GID>
<name>clear</name></connection>
<intersection>-55 1</intersection></vsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6.5,-16,6.5,-6</points>
<intersection>-16 8</intersection>
<intersection>-10.5 9</intersection>
<intersection>-9 2</intersection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6.5,-6,81.5,-6</points>
<intersection>6.5 0</intersection>
<intersection>31 7</intersection>
<intersection>56 3</intersection>
<intersection>81.5 6</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,-9,6.5,-9</points>
<connection>
<GID>92</GID>
<name>OUT_0</name></connection>
<intersection>6.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>56,-15,56,-6</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>-6 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>81.5,-14.5,81.5,-6</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>-6 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>31,-15.5,31,-6</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>-6 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>6.5,-16,7,-16</points>
<connection>
<GID>96</GID>
<name>IN_1</name></connection>
<intersection>6.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>6.5,-10.5,10,-10.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>6.5 0</intersection></hsegment></shape></wire></page 8>
<page 9>
<PageViewport>-9,45,113.4,-15.5</PageViewport>
<gate>
<ID>193</ID>
<type>AA_TOGGLE</type>
<position>1.5,1.5</position>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>207</ID>
<type>BB_CLOCK</type>
<position>0,21.5</position>
<output>
<ID>CLK</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_TOGGLE</type>
<position>1,-4</position>
<output>
<ID>OUT_0</ID>114 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>54,43</position>
<gparam>LABEL_TEXT UNIVERSAL SHIFT REGISTER</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>11,-12</position>
<gparam>LABEL_TEXT I3</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AE_MUX_4x1</type>
<position>17.5,2.5</position>
<input>
<ID>IN_0</ID>116 </input>
<input>
<ID>IN_1</ID>114 </input>
<input>
<ID>IN_2</ID>109 </input>
<input>
<ID>IN_3</ID>69 </input>
<output>
<ID>OUT</ID>122 </output>
<input>
<ID>SEL_0</ID>120 </input>
<input>
<ID>SEL_1</ID>126 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>101.5,-11</position>
<output>
<ID>OUT_0</ID>115 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>100</ID>
<type>AE_MUX_4x1</type>
<position>44,2.5</position>
<input>
<ID>IN_0</ID>117 </input>
<input>
<ID>IN_1</ID>116 </input>
<input>
<ID>IN_2</ID>118 </input>
<input>
<ID>IN_3</ID>97 </input>
<output>
<ID>OUT</ID>123 </output>
<input>
<ID>SEL_0</ID>120 </input>
<input>
<ID>SEL_1</ID>126 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>114</ID>
<type>AE_MUX_4x1</type>
<position>71,3.5</position>
<input>
<ID>IN_0</ID>118 </input>
<input>
<ID>IN_1</ID>117 </input>
<input>
<ID>IN_2</ID>113 </input>
<input>
<ID>IN_3</ID>98 </input>
<output>
<ID>OUT</ID>124 </output>
<input>
<ID>SEL_0</ID>120 </input>
<input>
<ID>SEL_1</ID>126 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>35,-10</position>
<gparam>LABEL_TEXT I2</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AE_MUX_4x1</type>
<position>100.5,3.5</position>
<input>
<ID>IN_0</ID>113 </input>
<input>
<ID>IN_1</ID>118 </input>
<input>
<ID>IN_2</ID>115 </input>
<input>
<ID>IN_3</ID>105 </input>
<output>
<ID>OUT</ID>125 </output>
<input>
<ID>SEL_0</ID>120 </input>
<input>
<ID>SEL_1</ID>126 </input>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>140</ID>
<type>AE_DFF_LOW</type>
<position>16.5,28.5</position>
<input>
<ID>IN_0</ID>122 </input>
<output>
<ID>OUT_0</ID>116 </output>
<input>
<ID>clear</ID>129 </input>
<input>
<ID>clock</ID>121 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_LABEL</type>
<position>64,-10.5</position>
<gparam>LABEL_TEXT I1</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>AA_LABEL</type>
<position>93.5,-11</position>
<gparam>LABEL_TEXT I0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>AE_DFF_LOW</type>
<position>42.5,28.5</position>
<input>
<ID>IN_0</ID>123 </input>
<output>
<ID>OUT_0</ID>109 </output>
<input>
<ID>clear</ID>129 </input>
<input>
<ID>clock</ID>121 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>158</ID>
<type>AE_DFF_LOW</type>
<position>71,28.5</position>
<input>
<ID>IN_0</ID>124 </input>
<output>
<ID>OUT_0</ID>118 </output>
<input>
<ID>clear</ID>129 </input>
<input>
<ID>clock</ID>121 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_LABEL</type>
<position>1.5,-7</position>
<gparam>LABEL_TEXT SERIAL INPUT</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>AE_DFF_LOW</type>
<position>99.5,28.5</position>
<input>
<ID>IN_0</ID>125 </input>
<output>
<ID>OUT_0</ID>119 </output>
<input>
<ID>clear</ID>129 </input>
<input>
<ID>clock</ID>121 </input>
<gparam>angle 90</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>164</ID>
<type>AA_TOGGLE</type>
<position>14.5,-10.5</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_LABEL</type>
<position>1,-9</position>
<gparam>LABEL_TEXT RIGHT SHIFT</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AA_TOGGLE</type>
<position>41,-11</position>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_TOGGLE</type>
<position>68,-11.5</position>
<output>
<ID>OUT_0</ID>98 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>0.5,18</position>
<gparam>LABEL_TEXT CLOCK PULSE</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>AA_TOGGLE</type>
<position>97.5,-12</position>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 90</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>175</ID>
<type>GA_LED</type>
<position>16,38</position>
<input>
<ID>N_in1</ID>116 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>AA_LABEL</type>
<position>-0.5,27</position>
<gparam>LABEL_TEXT CLEAR</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>GA_LED</type>
<position>42.5,38</position>
<input>
<ID>N_in1</ID>117 </input>
<input>
<ID>N_in2</ID>109 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>179</ID>
<type>GA_LED</type>
<position>70,37.5</position>
<input>
<ID>N_in1</ID>118 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>4,38</position>
<gparam>LABEL_TEXT PARALLEL OUTPUT BITS</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>181</ID>
<type>GA_LED</type>
<position>99.5,38</position>
<input>
<ID>N_in0</ID>119 </input>
<input>
<ID>N_in1</ID>113 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>AA_TOGGLE</type>
<position>-0.5,29.5</position>
<output>
<ID>OUT_0</ID>129 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>-1.5,6</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>-1.5,1.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>191</ID>
<type>AA_TOGGLE</type>
<position>2.5,6</position>
<output>
<ID>OUT_0</ID>120 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-8.5,14.5,-0.5</points>
<connection>
<GID>88</GID>
<name>IN_3</name></connection>
<connection>
<GID>164</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-9,41,-0.5</points>
<connection>
<GID>100</GID>
<name>IN_3</name></connection>
<connection>
<GID>168</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-9.5,68,0.5</points>
<connection>
<GID>114</GID>
<name>IN_3</name></connection>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-10,97.5,0.5</points>
<connection>
<GID>130</GID>
<name>IN_3</name></connection>
<connection>
<GID>173</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-2,36.5,38</points>
<intersection>-2 3</intersection>
<intersection>38 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>16.5,-2,36.5,-2</points>
<intersection>16.5 5</intersection>
<intersection>36.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>36.5,38,42.5,38</points>
<intersection>36.5 0</intersection>
<intersection>40.5 7</intersection>
<intersection>42.5 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>16.5,-2,16.5,-0.5</points>
<connection>
<GID>88</GID>
<name>IN_2</name></connection>
<intersection>-2 3</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>42.5,37,42.5,38</points>
<connection>
<GID>177</GID>
<name>N_in2</name></connection>
<intersection>38 4</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>40.5,31.5,40.5,38</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<intersection>38 4</intersection></vsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-6,90,15</points>
<intersection>-6 3</intersection>
<intersection>15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,15,108,15</points>
<intersection>90 0</intersection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>108,15,108,38</points>
<intersection>15 1</intersection>
<intersection>38 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>70,-6,103.5,-6</points>
<intersection>70 5</intersection>
<intersection>90 0</intersection>
<intersection>103.5 7</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>100.5,38,108,38</points>
<connection>
<GID>181</GID>
<name>N_in1</name></connection>
<intersection>108 2</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>70,-6,70,0.5</points>
<connection>
<GID>114</GID>
<name>IN_2</name></connection>
<intersection>-6 3</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>103.5,-6,103.5,0.5</points>
<connection>
<GID>130</GID>
<name>IN_0</name></connection>
<intersection>-6 3</intersection></vsegment></shape></wire>
<wire>
<ID>114</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18.5,-4,18.5,-0.5</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>3,-4,18.5,-4</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-4,99.5,0.5</points>
<connection>
<GID>130</GID>
<name>IN_2</name></connection>
<intersection>-4 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>101.5,-9,101.5,-4</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>99.5,-4,101.5,-4</points>
<intersection>99.5 0</intersection>
<intersection>101.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-3.5,26.5,38</points>
<intersection>-3.5 2</intersection>
<intersection>38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17,38,26.5,38</points>
<connection>
<GID>175</GID>
<name>N_in1</name></connection>
<intersection>19 3</intersection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20.5,-3.5,45,-3.5</points>
<intersection>20.5 7</intersection>
<intersection>26.5 0</intersection>
<intersection>45 6</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19,31.5,19,38</points>
<intersection>31.5 4</intersection>
<intersection>38 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>14.5,31.5,19,31.5</points>
<connection>
<GID>140</GID>
<name>OUT_0</name></connection>
<intersection>19 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>45,-3.5,45,-0.5</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>-3.5 2</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>20.5,-3.5,20.5,-0.5</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>-3.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-4,72,0.5</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>-4 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>51.5,-4,51.5,38</points>
<intersection>-4 2</intersection>
<intersection>38 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47,-4,72,-4</points>
<intersection>47 5</intersection>
<intersection>51.5 1</intersection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>43.5,38,51.5,38</points>
<connection>
<GID>177</GID>
<name>N_in1</name></connection>
<intersection>51.5 1</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>47,-4,47,-0.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>-4 2</intersection></vsegment></shape></wire>
<wire>
<ID>118</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>74,-2.5,101.5,-2.5</points>
<intersection>74 12</intersection>
<intersection>83 3</intersection>
<intersection>101.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>83,-2.5,83,37.5</points>
<intersection>-2.5 2</intersection>
<intersection>37.5 5</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>101.5,-2.5,101.5,0.5</points>
<connection>
<GID>130</GID>
<name>IN_1</name></connection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>61,37.5,83,37.5</points>
<connection>
<GID>179</GID>
<name>N_in1</name></connection>
<intersection>61 8</intersection>
<intersection>69 10</intersection>
<intersection>83 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>43,-6,43,-0.5</points>
<connection>
<GID>100</GID>
<name>IN_2</name></connection>
<intersection>-6 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>43,-6,61,-6</points>
<intersection>43 6</intersection>
<intersection>61 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>61,-6,61,37.5</points>
<intersection>-6 7</intersection>
<intersection>37.5 5</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>69,31.5,69,37.5</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<intersection>37.5 5</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>74,-2.5,74,0.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>-2.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>93.5,31.5,93.5,38</points>
<intersection>31.5 2</intersection>
<intersection>38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>93.5,38,98.5,38</points>
<connection>
<GID>181</GID>
<name>N_in0</name></connection>
<intersection>93.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93.5,31.5,97.5,31.5</points>
<connection>
<GID>162</GID>
<name>OUT_0</name></connection>
<intersection>93.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,6,8.5,9.5</points>
<intersection>6 2</intersection>
<intersection>9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,9.5,95.5,9.5</points>
<intersection>8.5 0</intersection>
<intersection>12.5 6</intersection>
<intersection>39 5</intersection>
<intersection>66 8</intersection>
<intersection>95.5 7</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4.5,6,8.5,6</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<intersection>8.5 0</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>39,3.5,39,9.5</points>
<connection>
<GID>100</GID>
<name>SEL_0</name></connection>
<intersection>9.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>12.5,3.5,12.5,9.5</points>
<connection>
<GID>88</GID>
<name>SEL_0</name></connection>
<intersection>9.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>95.5,4.5,95.5,9.5</points>
<connection>
<GID>130</GID>
<name>SEL_0</name></connection>
<intersection>9.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>66,4.5,66,9.5</points>
<connection>
<GID>114</GID>
<name>SEL_0</name></connection>
<intersection>9.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,21.5,17.5,25.5</points>
<connection>
<GID>140</GID>
<name>clock</name></connection>
<intersection>21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>4,21.5,100.5,21.5</points>
<connection>
<GID>207</GID>
<name>CLK</name></connection>
<intersection>17.5 0</intersection>
<intersection>43.5 3</intersection>
<intersection>72 5</intersection>
<intersection>100.5 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43.5,21.5,43.5,25.5</points>
<connection>
<GID>154</GID>
<name>clock</name></connection>
<intersection>21.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>72,21.5,72,25.5</points>
<connection>
<GID>158</GID>
<name>clock</name></connection>
<intersection>21.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>100.5,21.5,100.5,25.5</points>
<connection>
<GID>162</GID>
<name>clock</name></connection>
<intersection>21.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,15.5,14.5,25.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>15.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>17.5,5.5,17.5,15.5</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<intersection>15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>14.5,15.5,17.5,15.5</points>
<intersection>14.5 0</intersection>
<intersection>17.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>123</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,15.5,40.5,25.5</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>15.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>44,5.5,44,15.5</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<intersection>15.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>40.5,15.5,44,15.5</points>
<intersection>40.5 0</intersection>
<intersection>44 1</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,16,69,25.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>16 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>71,6.5,71,16</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>69,16,71,16</points>
<intersection>69 0</intersection>
<intersection>71 1</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,16,97.5,25.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>16 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>100.5,6.5,100.5,16</points>
<connection>
<GID>130</GID>
<name>OUT</name></connection>
<intersection>16 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>97.5,16,100.5,16</points>
<intersection>97.5 0</intersection>
<intersection>100.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,1.5,8,6</points>
<intersection>1.5 2</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,6,94.5,6</points>
<intersection>8 0</intersection>
<intersection>12.5 7</intersection>
<intersection>39 6</intersection>
<intersection>66 4</intersection>
<intersection>94.5 8</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>3.5,1.5,8,1.5</points>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection>
<intersection>8 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>66,3.5,66,6</points>
<connection>
<GID>114</GID>
<name>SEL_1</name></connection>
<intersection>6 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>39,2.5,39,6</points>
<connection>
<GID>100</GID>
<name>SEL_1</name></connection>
<intersection>6 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>12.5,2.5,12.5,6</points>
<connection>
<GID>88</GID>
<name>SEL_1</name></connection>
<intersection>6 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>94.5,3.5,94.5,6</points>
<intersection>3.5 9</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>94.5,3.5,95.5,3.5</points>
<connection>
<GID>130</GID>
<name>SEL_1</name></connection>
<intersection>94.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1.5,33.5,105.5,33.5</points>
<intersection>1.5 12</intersection>
<intersection>23.5 3</intersection>
<intersection>48.5 6</intersection>
<intersection>75 8</intersection>
<intersection>105.5 10</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>23.5,28.5,23.5,33.5</points>
<intersection>28.5 13</intersection>
<intersection>33.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>48.5,28.5,48.5,33.5</points>
<intersection>28.5 14</intersection>
<intersection>33.5 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>75,28.5,75,33.5</points>
<connection>
<GID>158</GID>
<name>clear</name></connection>
<intersection>33.5 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>105.5,28.5,105.5,33.5</points>
<intersection>28.5 15</intersection>
<intersection>33.5 1</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>1.5,29.5,1.5,33.5</points>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection>
<intersection>33.5 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>20.5,28.5,23.5,28.5</points>
<connection>
<GID>140</GID>
<name>clear</name></connection>
<intersection>23.5 3</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>46.5,28.5,48.5,28.5</points>
<connection>
<GID>154</GID>
<name>clear</name></connection>
<intersection>48.5 6</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>103.5,28.5,105.5,28.5</points>
<connection>
<GID>162</GID>
<name>clear</name></connection>
<intersection>105.5 10</intersection></hsegment></shape></wire></page 9></circuit>