<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>1187.51,1515.9,1405.73,1408.04</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>1229.5,1503.5</position>
<gparam>LABEL_TEXT HALF ADDER</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AI_XOR2</type>
<position>1227,1473.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>1344.5,1504</position>
<gparam>LABEL_TEXT HALF SUBTRACTOR</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>1367,1479.5</position>
<gparam>LABEL_TEXT DIFFERENCE</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>1367.5,1456.5</position>
<gparam>LABEL_TEXT BORROW</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>1217,1439</position>
<gparam>LABEL_TEXT SUM=X'Y+XY'</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>1217.5,1432</position>
<gparam>LABEL_TEXT SUM=X(XOR)Y</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_LABEL</type>
<position>1217,1424.5</position>
<gparam>LABEL_TEXT CARRY=XY</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>1329,1440.5</position>
<gparam>LABEL_TEXT DIFFERENCE=X'Y+XY'</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>1328.5,1432.5</position>
<gparam>LABEL_TEXT DIFFERENCE=X(XOR)Y</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>1329.5,1423</position>
<gparam>LABEL_TEXT BORROW=X'Y</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>1228,1482</position>
<gparam>LABEL_TEXT SUM</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>1242.5,1450</position>
<gparam>LABEL_TEXT CARRY</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>1204.5,1482.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_AND2</type>
<position>1228,1456</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>1206,1467.5</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>GA_LED</type>
<position>1240.5,1474</position>
<input>
<ID>N_in0</ID>10 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>GA_LED</type>
<position>1241,1456.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>1197,1482.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>1209,1464</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AI_XOR2</type>
<position>1325.5,1478.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>1293,1485</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>1292,1474.5</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>1282.5,1486</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>1282.5,1476</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>GA_LED</type>
<position>1343,1478.5</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND2</type>
<position>1327.5,1456</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>GA_LED</type>
<position>1344,1456</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_INVERTER</type>
<position>1317,1468.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1308.5,1479.5,1308.5,1485</points>
<intersection>1479.5 1</intersection>
<intersection>1485 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1308.5,1479.5,1322.5,1479.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>1308.5 0</intersection>
<intersection>1314 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1295,1485,1308.5,1485</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>1308.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1314,1468.5,1314,1479.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>1479.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1322,1457,1322,1468.5</points>
<intersection>1457 1</intersection>
<intersection>1468.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1322,1457,1324.5,1457</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>1322 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1320,1468.5,1322,1468.5</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>1322 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1215,1474.5,1215,1482.5</points>
<intersection>1474.5 1</intersection>
<intersection>1482.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1200,1474.5,1224,1474.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>1200 3</intersection>
<intersection>1215 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1206.5,1482.5,1215,1482.5</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>1215 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1200,1457,1200,1474.5</points>
<intersection>1457 4</intersection>
<intersection>1474.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1200,1457,1225,1457</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>1200 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1216,1455,1216,1472.5</points>
<intersection>1455 3</intersection>
<intersection>1467.5 2</intersection>
<intersection>1472.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1216,1472.5,1224,1472.5</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>1216 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1208,1467.5,1216,1467.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>1216 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>1216,1455,1225,1455</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>1216 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1231,1456,1240,1456</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>1240 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1240,1456,1240,1456.5</points>
<connection>
<GID>32</GID>
<name>N_in0</name></connection>
<intersection>1456 1</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1230,1473.5,1239.5,1473.5</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>1239.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1239.5,1473.5,1239.5,1474</points>
<connection>
<GID>30</GID>
<name>N_in0</name></connection>
<intersection>1473.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>1308,1474.5,1308,1477.5</points>
<intersection>1474.5 2</intersection>
<intersection>1477.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1308,1477.5,1322.5,1477.5</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>1308 0</intersection>
<intersection>1310.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>1294,1474.5,1308,1474.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>1308 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>1310.5,1449.5,1310.5,1477.5</points>
<intersection>1449.5 4</intersection>
<intersection>1477.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>1310.5,1449.5,1324.5,1449.5</points>
<intersection>1310.5 3</intersection>
<intersection>1324.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>1324.5,1449.5,1324.5,1455</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>1449.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1328.5,1478.5,1342,1478.5</points>
<connection>
<GID>48</GID>
<name>N_in0</name></connection>
<connection>
<GID>38</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>1330.5,1456,1343,1456</points>
<connection>
<GID>54</GID>
<name>N_in0</name></connection>
<connection>
<GID>50</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>74.2142,22.1877,217.447,-48.6096</PageViewport>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>206.5,-16</position>
<gparam>LABEL_TEXT CARRY</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>136,-31.5</position>
<gparam>LABEL_TEXT SUM=X(XOR)Y(XOR)Z</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>138,-39</position>
<gparam>LABEL_TEXT CARRY=X(XOR)Y(XOR)Z+XY</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>109.5,-6</position>
<gparam>LABEL_TEXT XY</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>138,-20.5</position>
<gparam>LABEL_TEXT X(XOR)Y(XOR)Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>139,16.5</position>
<gparam>LABEL_TEXT FULL ADDER</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AI_XOR2</type>
<position>110,0</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_LABEL</type>
<position>177,-12</position>
<gparam>LABEL_TEXT X(XOR)Y(XOR)Z+XY</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AI_XOR2</type>
<position>153,0</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_TOGGLE</type>
<position>88,5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_TOGGLE</type>
<position>88,-2.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>82,5.5</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>82,-2</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AA_TOGGLE</type>
<position>88.5,-17.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>83,-16.5</position>
<gparam>LABEL_TEXT Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>199.5,0</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>206,0.5</position>
<gparam>LABEL_TEXT SUM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>110,6.5</position>
<gparam>LABEL_TEXT X(XOR)Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>174,4</position>
<gparam>LABEL_TEXT X(XOR)Y(XOR)Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_AND2</type>
<position>108.5,-11</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_AND2</type>
<position>140,-16.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>AE_OR2</type>
<position>158,-16.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>GA_LED</type>
<position>198.5,-16.5</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,1,98.5,5</points>
<intersection>1 1</intersection>
<intersection>5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,1,107,1</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>98.5 0</intersection>
<intersection>101 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90,5,98.5,5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>101,-10,101,1</points>
<intersection>-10 4</intersection>
<intersection>1 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>101,-10,105.5,-10</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>101 3</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,-2.5,107,-2.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<intersection>93 6</intersection>
<intersection>107 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>107,-2.5,107,-1</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>93,-12,93,-2.5</points>
<intersection>-12 7</intersection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>93,-12,105.5,-12</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<intersection>93 6</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-15.5,129.5,4.5</points>
<intersection>-15.5 5</intersection>
<intersection>0 2</intersection>
<intersection>4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,4.5,146,4.5</points>
<intersection>129.5 0</intersection>
<intersection>146 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>113,0,129.5,0</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>129.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>146,1,146,4.5</points>
<intersection>1 4</intersection>
<intersection>4.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>146,1,150,1</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>146 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>129.5,-15.5,137,-15.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120,-17.5,120,-7.5</points>
<intersection>-17.5 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>120,-7.5,146,-7.5</points>
<intersection>120 0</intersection>
<intersection>146 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-17.5,137,-17.5</points>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>120 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>146,-7.5,146,-1</points>
<intersection>-7.5 1</intersection>
<intersection>-1 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>146,-1,150,-1</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>146 3</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>156,0,198.5,0</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<connection>
<GID>59</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,-17.5,149,-16.5</points>
<intersection>-17.5 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149,-17.5,155,-17.5</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>149 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>143,-16.5,149,-16.5</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>149 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>111.5,-11,155,-11</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>155 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>155,-15.5,155,-11</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>-11 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>161,-16.5,197.5,-16.5</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<connection>
<GID>75</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>122.874,44.9149,266.107,-25.8824</PageViewport>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>191,40</position>
<gparam>LABEL_TEXT FULL SUBTRACTOR</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AI_XOR2</type>
<position>161,23</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AI_XOR2</type>
<position>203.5,23.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>138,32</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_TOGGLE</type>
<position>138.5,19.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>138.5,-0.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>134,31</position>
<gparam>LABEL_TEXT X</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>134.5,20.5</position>
<gparam>LABEL_TEXT Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>151,30.5</position>
<gparam>LABEL_TEXT X(XOR)Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>133,0</position>
<gparam>LABEL_TEXT Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>GA_LED</type>
<position>240,23.5</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>221,27</position>
<gparam>LABEL_TEXT X(XOR)Y(XOR)Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>253,24.5</position>
<gparam>LABEL_TEXT DIFFERENCE</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_AND2</type>
<position>159.5,10.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>87</ID>
<type>AA_INVERTER</type>
<position>143,11.5</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>158,5</position>
<gparam>LABEL_TEXT Z(XOR)(X+Y)'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_AND2</type>
<position>200.5,-7</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>AE_OR2</type>
<position>218,9.5</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_INVERTER</type>
<position>168,-4</position>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>97</ID>
<type>GA_LED</type>
<position>241,10.5</position>
<input>
<ID>N_in0</ID>32 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>250.5,11</position>
<gparam>LABEL_TEXT BORROW</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>AA_LABEL</type>
<position>199.5,-1</position>
<gparam>LABEL_TEXT X'Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>AA_LABEL</type>
<position>230.5,5</position>
<gparam>LABEL_TEXT Z(X XOR Y)+XY'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>191,-13.5</position>
<gparam>LABEL_TEXT DIFFERENCE=X(XOR)Y(XOR)Z</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>193,-20.5</position>
<gparam>LABEL_TEXT BORROW=Z(X XOR Y)'+X'Y</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,19.5,149,22</points>
<intersection>19.5 2</intersection>
<intersection>22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>128.5,22,158,22</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>128.5 3</intersection>
<intersection>149 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140.5,19.5,149,19.5</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<intersection>149 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>128.5,-8,128.5,22</points>
<intersection>-8 4</intersection>
<intersection>22 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>128.5,-8,197.5,-8</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>128.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-0.5,170.5,6</points>
<intersection>-0.5 2</intersection>
<intersection>6 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170.5,6,197,6</points>
<intersection>170.5 0</intersection>
<intersection>197 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140.5,-0.5,170.5,-0.5</points>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection>
<intersection>145.5 5</intersection>
<intersection>170.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>197,6,197,22.5</points>
<intersection>6 1</intersection>
<intersection>22.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>197,22.5,200.5,22.5</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>197 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>145.5,-0.5,145.5,9.5</points>
<intersection>-0.5 2</intersection>
<intersection>9.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>145.5,9.5,156.5,9.5</points>
<connection>
<GID>85</GID>
<name>IN_1</name></connection>
<intersection>145.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>206.5,23.5,239,23.5</points>
<connection>
<GID>79</GID>
<name>N_in0</name></connection>
<connection>
<GID>52</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>146,11.5,156.5,11.5</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>162.5,10.5,215,10.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<connection>
<GID>85</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>182,16,182,24.5</points>
<intersection>16 2</intersection>
<intersection>24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>182,24.5,200.5,24.5</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>182 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140,16,182,16</points>
<intersection>140 3</intersection>
<intersection>164 4</intersection>
<intersection>182 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>140,11.5,140,16</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>16 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>164,16,164,23</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>16 2</intersection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>126,-4,126,25.5</points>
<intersection>-4 2</intersection>
<intersection>25.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>126,25.5,155,25.5</points>
<intersection>126 0</intersection>
<intersection>141 3</intersection>
<intersection>155 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>126,-4,165,-4</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>126 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>141,25.5,141,32</points>
<intersection>25.5 1</intersection>
<intersection>32 6</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>155,24,155,25.5</points>
<intersection>24 5</intersection>
<intersection>25.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>155,24,158,24</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>155 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>140,32,141,32</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>141 3</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>184,-6,184,-4</points>
<intersection>-6 1</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>184,-6,197.5,-6</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>184 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>171,-4,184,-4</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<intersection>184 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>209,-7,209,8.5</points>
<intersection>-7 2</intersection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>209,8.5,215,8.5</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>209 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>203.5,-7,209,-7</points>
<connection>
<GID>91</GID>
<name>OUT</name></connection>
<intersection>209 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>221,9.5,240,9.5</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<intersection>240 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>240,9.5,240,10.5</points>
<connection>
<GID>97</GID>
<name>N_in0</name></connection>
<intersection>9.5 1</intersection></vsegment></shape></wire></page 2>
<page 3>
<PageViewport>18.0222,43.5464,161.255,-27.2509</PageViewport></page 3>
<page 4>
<PageViewport>-0.280104,33.7194,339.234,-134.096</PageViewport></page 4>
<page 5>
<PageViewport>-0.280104,33.7194,339.234,-134.096</PageViewport></page 5>
<page 6>
<PageViewport>-0.280104,33.7194,339.234,-134.096</PageViewport></page 6>
<page 7>
<PageViewport>-0.280104,33.7194,339.234,-134.096</PageViewport></page 7>
<page 8>
<PageViewport>-0.280104,33.7194,339.234,-134.096</PageViewport></page 8>
<page 9>
<PageViewport>-0.280104,33.7194,339.234,-134.096</PageViewport></page 9></circuit>