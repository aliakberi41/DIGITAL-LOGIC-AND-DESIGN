<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>0,3,122.4,-57.5</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>22,-1.5</position>
<gparam>LABEL_TEXT HALF ADDER</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>GA_LED</type>
<position>34.5,-19.5</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>90.5,-2</position>
<gparam>LABEL_TEXT HALF SUBTRACTOR</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AI_XOR2</type>
<position>22,-20.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>GA_LED</type>
<position>35,-32</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_TOGGLE</type>
<position>9,-13</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>6,-25.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>11</ID>
<type>GA_LED</type>
<position>103,-19</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>24,-32.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AI_XOR2</type>
<position>85.5,-19</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>GA_LED</type>
<position>104,-34.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>92.5,-35</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>65,-13</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>64.5,-23</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_INVERTER</type>
<position>83,-28.5</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>19,-41.5</position>
<gparam>LABEL_TEXT SUM=X(XOR)Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>18.5,-47</position>
<gparam>LABEL_TEXT CARRY=XY</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>87,-41</position>
<gparam>LABEL_TEXT DIFFERENCE=X(XOR)Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>88,-46</position>
<gparam>LABEL_TEXT BORROW=X'Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-19.5,15,-13</points>
<intersection>-19.5 1</intersection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15,-19.5,19,-19.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection>
<intersection>17 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-13,15,-13</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>15 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>17,-31.5,17,-19.5</points>
<intersection>-31.5 4</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>17,-31.5,21,-31.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>17 3</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-33.5,14.5,-21.5</points>
<intersection>-33.5 3</intersection>
<intersection>-25.5 2</intersection>
<intersection>-21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-21.5,19,-21.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8,-25.5,14.5,-25.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>14.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>14.5,-33.5,21,-33.5</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-18,74.5,-13</points>
<intersection>-18 1</intersection>
<intersection>-13 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-18,82.5,-18</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>74.5 0</intersection>
<intersection>80 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>67,-13,74.5,-13</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>80,-28.5,80,-18</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>-18 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-23,74.5,-20</points>
<intersection>-23 2</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-20,82.5,-20</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection>
<intersection>76.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66.5,-23,74.5,-23</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>74.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>76.5,-36,76.5,-20</points>
<intersection>-36 4</intersection>
<intersection>-20 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>76.5,-36,89.5,-36</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>76.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86,-34,86,-28.5</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86,-34,89.5,-34</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>86 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30.5,-32.5,30.5,-32</points>
<intersection>-32.5 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-32,34,-32</points>
<connection>
<GID>7</GID>
<name>N_in0</name></connection>
<intersection>30.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,-32.5,30.5,-32.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>30.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-20.5,29,-19.5</points>
<intersection>-20.5 2</intersection>
<intersection>-19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-19.5,33.5,-19.5</points>
<connection>
<GID>3</GID>
<name>N_in0</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-20.5,29,-20.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88.5,-19,102,-19</points>
<connection>
<GID>11</GID>
<name>N_in0</name></connection>
<connection>
<GID>14</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99,-35,99,-34.5</points>
<intersection>-35 2</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99,-34.5,103,-34.5</points>
<connection>
<GID>15</GID>
<name>N_in0</name></connection>
<intersection>99 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,-35,99,-35</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>99 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>88.5,-16.5</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>GA_LED</type>
<position>92.5,-32</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>AA_LABEL</type>
<position>73.5,-47</position>
<gparam>LABEL_TEXT SUM=X(XOR)Y(XOR)Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>73.5,-51.5</position>
<gparam>LABEL_TEXT CARRY=X(XOR)Y(XOR)Z+XY</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>55,-4</position>
<gparam>LABEL_TEXT FULL ADDERS</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AI_XOR2</type>
<position>29.5,-18</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AI_XOR2</type>
<position>72,-17.5</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_TOGGLE</type>
<position>6.5,-10.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>6.5,-20.5</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>6.5,-44.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>28,-31.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_AND2</type>
<position>67.5,-32</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AE_OR2</type>
<position>82.5,-32</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-17,17.5,-10.5</points>
<intersection>-17 1</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-17,26.5,-17</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection>
<intersection>22 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-10.5,17.5,-10.5</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22,-30.5,22,-17</points>
<intersection>-30.5 4</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>22,-30.5,25,-30.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>22 3</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-20.5,17.5,-19</points>
<intersection>-20.5 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>17.5,-19,26.5,-19</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>17.5 0</intersection>
<intersection>20 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-20.5,17.5,-20.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20,-32.5,20,-19</points>
<intersection>-32.5 4</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20,-32.5,25,-32.5</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>20 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-12.5,60.5,-12.5</points>
<intersection>35.5 4</intersection>
<intersection>60.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>60.5,-31,60.5,-12.5</points>
<intersection>-31 6</intersection>
<intersection>-16.5 7</intersection>
<intersection>-12.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>35.5,-18,35.5,-12.5</points>
<intersection>-18 5</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>32.5,-18,35.5,-18</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>35.5 4</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>60.5,-31,64.5,-31</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>60.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>60.5,-16.5,69,-16.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>60.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-44.5,50.5,-18.5</points>
<intersection>-44.5 2</intersection>
<intersection>-33 5</intersection>
<intersection>-18.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-44.5,50.5,-44.5</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>50.5,-18.5,69,-18.5</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>50.5,-33,64.5,-33</points>
<connection>
<GID>46</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-32,75,-31</points>
<intersection>-32 2</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-31,79.5,-31</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-32,75,-32</points>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-39,79.5,-39</points>
<intersection>31 3</intersection>
<intersection>79.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>31,-39,31,-31.5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>-39 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>79.5,-39,79.5,-33</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>-39 1</intersection></vsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-17.5,81,-16.5</points>
<intersection>-17.5 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,-16.5,87.5,-16.5</points>
<connection>
<GID>19</GID>
<name>N_in0</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>75,-17.5,81,-17.5</points>
<connection>
<GID>36</GID>
<name>OUT</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>85.5,-32,91.5,-32</points>
<connection>
<GID>23</GID>
<name>N_in0</name></connection>
<connection>
<GID>48</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport>
<gate>
<ID>5</ID>
<type>GA_LED</type>
<position>89.5,-18.5</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>81.5,-47</position>
<gparam>LABEL_TEXT DIFFERENCE=X(XOR)(Y(XOR)Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_AND2</type>
<position>65,-35</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_INVERTER</type>
<position>45,-27.5</position>
<input>
<ID>IN_0</ID>20 </input>
<output>
<ID>OUT_0</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>82,-51.5</position>
<gparam>LABEL_TEXT BORROW=(X+Y)'XOR(Z)+X'Y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AE_OR2</type>
<position>79.5,-35.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>56.5,-4</position>
<gparam>LABEL_TEXT FULL SUBTRACTORS</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>GA_LED</type>
<position>90,-35</position>
<input>
<ID>N_in0</ID>27 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AI_XOR2</type>
<position>31,-19.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>43</ID>
<type>AI_XOR2</type>
<position>70,-19</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AA_TOGGLE</type>
<position>10,-11.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>10,-24.5</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_TOGGLE</type>
<position>10.5,-49</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_INVERTER</type>
<position>28.5,-28.5</position>
<input>
<ID>IN_0</ID>18 </input>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_AND2</type>
<position>37,-35.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>19 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-18.5,20,-11.5</points>
<intersection>-18.5 1</intersection>
<intersection>-11.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-18.5,28,-18.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>20 0</intersection>
<intersection>25.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-11.5,20,-11.5</points>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>20 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25.5,-28.5,25.5,-18.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>-18.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20,-24.5,20,-20.5</points>
<intersection>-24.5 2</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20,-20.5,28,-20.5</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>20 0</intersection>
<intersection>22.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-24.5,20,-24.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>20 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22.5,-36.5,22.5,-20.5</points>
<intersection>-36.5 4</intersection>
<intersection>-20.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>22.5,-36.5,34,-36.5</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>22.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-19.5,50.5,-18</points>
<intersection>-19.5 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-18,67,-18</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-19.5,50.5,-19.5</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>42 3</intersection>
<intersection>50.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>42,-27.5,42,-19.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-19.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-49,52.5,-20</points>
<intersection>-49 2</intersection>
<intersection>-36 5</intersection>
<intersection>-20 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-49,52.5,-49</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>52.5,-20,67,-20</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>52.5,-36,62,-36</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-34.5,33,-28.5</points>
<intersection>-34.5 1</intersection>
<intersection>-28.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-34.5,34,-34.5</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31.5,-28.5,33,-28.5</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-19,80.5,-18.5</points>
<intersection>-19 2</intersection>
<intersection>-18.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-18.5,88.5,-18.5</points>
<connection>
<GID>5</GID>
<name>N_in0</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73,-19,80.5,-19</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-34,55,-27.5</points>
<intersection>-34 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-34,62,-34</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-27.5,55,-27.5</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72,-35,72,-34.5</points>
<intersection>-35 2</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72,-34.5,76.5,-34.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>72 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-35,72,-35</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>72 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>40,-41,76.5,-41</points>
<intersection>40 3</intersection>
<intersection>76.5 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>40,-41,40,-35.5</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>-41 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>76.5,-41,76.5,-36.5</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>-41 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85.5,-35.5,85.5,-35</points>
<intersection>-35.5 2</intersection>
<intersection>-35 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-35,89,-35</points>
<connection>
<GID>37</GID>
<name>N_in0</name></connection>
<intersection>85.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-35.5,85.5,-35.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>85.5 0</intersection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-23.4,16.0667,139.8,-64.6</PageViewport>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>79.5,-9</position>
<gparam>LABEL_TEXT D0=X'Y'Z'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>44.5,12</position>
<gparam>LABEL_TEXT DECODERS</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>79,-15</position>
<gparam>LABEL_TEXT D1=X'Y'Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>79.5,-21.5</position>
<gparam>LABEL_TEXT D2=X'YZ'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>79,-27.5</position>
<gparam>LABEL_TEXT D3=X'YZ</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>-9.5,0</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_TOGGLE</type>
<position>-9.5,-16</position>
<output>
<ID>OUT_0</ID>51 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>79.5,-33</position>
<gparam>LABEL_TEXT D4=XY'Z'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_TOGGLE</type>
<position>-9.5,-35</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>79,-39.5</position>
<gparam>LABEL_TEXT D5=XY'Z</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>79.5,-45.5</position>
<gparam>LABEL_TEXT D6=XYZ'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>79,-53.5</position>
<gparam>LABEL_TEXT D7=XYZ</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>72,11.5</position>
<gparam>LABEL_TEXT (3*8)</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>GA_LED</type>
<position>65.5,-10</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>65.5,-16</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>GA_LED</type>
<position>65.5,-21.5</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>GA_LED</type>
<position>65.5,-27.5</position>
<input>
<ID>N_in0</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>GA_LED</type>
<position>65.5,-33.5</position>
<input>
<ID>N_in0</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>GA_LED</type>
<position>65.5,-40</position>
<input>
<ID>N_in0</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>GA_LED</type>
<position>65.5,-46.5</position>
<input>
<ID>N_in0</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>GA_LED</type>
<position>66,-54.5</position>
<input>
<ID>N_in0</ID>49 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>95</ID>
<type>AA_AND3</type>
<position>32.5,2</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>56 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_AND3</type>
<position>32.5,-7</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>52 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_AND3</type>
<position>32.5,-16</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>56 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_AND3</type>
<position>32.5,-23.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>52 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_AND3</type>
<position>32.5,-32</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>56 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>105</ID>
<type>AA_AND3</type>
<position>32.5,-40</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>55 </input>
<input>
<ID>IN_2</ID>52 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>107</ID>
<type>AA_AND3</type>
<position>32.5,-48.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>56 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_AND3</type>
<position>32.5,-57.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>52 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_INVERTER</type>
<position>1,0.5</position>
<input>
<ID>IN_0</ID>50 </input>
<output>
<ID>OUT_0</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_INVERTER</type>
<position>1.5,-15.5</position>
<input>
<ID>IN_0</ID>51 </input>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_INVERTER</type>
<position>2,-35</position>
<input>
<ID>IN_0</ID>52 </input>
<output>
<ID>OUT_0</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-10,49.5,2</points>
<intersection>-10 1</intersection>
<intersection>2 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-10,64.5,-10</points>
<connection>
<GID>79</GID>
<name>N_in0</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,2,49.5,2</points>
<connection>
<GID>95</GID>
<name>OUT</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>48,-16,48,-7</points>
<intersection>-16 1</intersection>
<intersection>-7 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>48,-16,64.5,-16</points>
<connection>
<GID>81</GID>
<name>N_in0</name></connection>
<intersection>48 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-7,48,-7</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<intersection>48 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-21.5,45,-16</points>
<intersection>-21.5 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-21.5,64.5,-21.5</points>
<connection>
<GID>83</GID>
<name>N_in0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-16,45,-16</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-27.5,50,-23.5</points>
<intersection>-27.5 1</intersection>
<intersection>-23.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-27.5,64.5,-27.5</points>
<connection>
<GID>85</GID>
<name>N_in0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-23.5,50,-23.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-33.5,50,-32</points>
<intersection>-33.5 1</intersection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-33.5,64.5,-33.5</points>
<connection>
<GID>87</GID>
<name>N_in0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-32,50,-32</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-40,64.5,-40</points>
<connection>
<GID>89</GID>
<name>N_in0</name></connection>
<connection>
<GID>105</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-48.5,50,-46.5</points>
<intersection>-48.5 2</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-46.5,64.5,-46.5</points>
<connection>
<GID>91</GID>
<name>N_in0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-48.5,50,-48.5</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50,-57.5,50,-54.5</points>
<intersection>-57.5 2</intersection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-54.5,65,-54.5</points>
<connection>
<GID>93</GID>
<name>N_in0</name></connection>
<intersection>50 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-57.5,50,-57.5</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<intersection>50 0</intersection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,0,-4.5,7.5</points>
<intersection>0 2</intersection>
<intersection>7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,7.5,15.5,7.5</points>
<intersection>-4.5 0</intersection>
<intersection>-2 5</intersection>
<intersection>15.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,0,-4.5,0</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15.5,-55.5,15.5,7.5</points>
<intersection>-55.5 4</intersection>
<intersection>-30 6</intersection>
<intersection>7.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>15.5,-55.5,29.5,-55.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-2,0.5,-2,7.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>7.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>15.5,-30,29.5,-30</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection>
<intersection>26 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>26,-46.5,26,-30</points>
<intersection>-46.5 10</intersection>
<intersection>-38 8</intersection>
<intersection>-30 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>26,-38,29.5,-38</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>26 7</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>26,-46.5,29.5,-46.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>26 7</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-16,-4.5,-11</points>
<intersection>-16 2</intersection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4.5,-11,22.5,-11</points>
<intersection>-4.5 0</intersection>
<intersection>-1.5 4</intersection>
<intersection>22.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-16,-4.5,-16</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22.5,-57.5,22.5,-11</points>
<intersection>-57.5 9</intersection>
<intersection>-48.5 10</intersection>
<intersection>-23.5 6</intersection>
<intersection>-16 7</intersection>
<intersection>-11 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-1.5,-15.5,-1.5,-11</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>-11 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>22.5,-23.5,29.5,-23.5</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>22.5 3</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>22.5,-16,29.5,-16</points>
<connection>
<GID>99</GID>
<name>IN_1</name></connection>
<intersection>22.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>22.5,-57.5,29.5,-57.5</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<intersection>22.5 3</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>22.5,-48.5,29.5,-48.5</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>22.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-7.5,-25.5,29.5,-25.5</points>
<connection>
<GID>101</GID>
<name>IN_2</name></connection>
<intersection>-7.5 5</intersection>
<intersection>-1 4</intersection>
<intersection>13 2</intersection>
<intersection>19 7</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>13,-25.5,13,-9</points>
<intersection>-25.5 1</intersection>
<intersection>-9 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>13,-9,29.5,-9</points>
<connection>
<GID>97</GID>
<name>IN_2</name></connection>
<intersection>13 2</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-1,-35,-1,-25.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>-25.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-7.5,-35,-7.5,-25.5</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>-25.5 1</intersection></vsegment>
<vsegment>
<ID>7</ID>
<points>19,-59.5,19,-25.5</points>
<intersection>-59.5 10</intersection>
<intersection>-42 11</intersection>
<intersection>-25.5 1</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>19,-59.5,29.5,-59.5</points>
<connection>
<GID>109</GID>
<name>IN_2</name></connection>
<intersection>19 7</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>19,-42,29.5,-42</points>
<connection>
<GID>105</GID>
<name>IN_2</name></connection>
<intersection>19 7</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>4,4,29.5,4</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>4 3</intersection>
<intersection>24 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>4,0.5,4,4</points>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<intersection>4 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>24,-21.5,24,4</points>
<intersection>-21.5 9</intersection>
<intersection>-14 7</intersection>
<intersection>-5 5</intersection>
<intersection>4 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>24,-5,29.5,-5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<intersection>24 4</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>24,-14,29.5,-14</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<intersection>24 4</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>24,-21.5,29.5,-21.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>24 4</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>6,-15.5,6,2</points>
<intersection>-15.5 2</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>6,2,29.5,2</points>
<connection>
<GID>95</GID>
<name>IN_1</name></connection>
<intersection>6 0</intersection>
<intersection>20 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>4.5,-15.5,6,-15.5</points>
<connection>
<GID>113</GID>
<name>OUT_0</name></connection>
<intersection>6 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20,-7,20,2</points>
<intersection>-7 4</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20,-7,29.5,-7</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<intersection>20 3</intersection>
<intersection>26 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>26,-32,26,-7</points>
<intersection>-32 6</intersection>
<intersection>-7 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>24,-32,29.5,-32</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<intersection>24 7</intersection>
<intersection>26 5</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>24,-40,24,-32</points>
<intersection>-40 8</intersection>
<intersection>-32 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>24,-40,29.5,-40</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>24 7</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8,-35,8,0</points>
<intersection>-35 2</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,0,29.5,0</points>
<connection>
<GID>95</GID>
<name>IN_2</name></connection>
<intersection>8 0</intersection>
<intersection>17 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>5,-35,8,-35</points>
<connection>
<GID>115</GID>
<name>OUT_0</name></connection>
<intersection>8 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>17,-34,17,0</points>
<intersection>-34 6</intersection>
<intersection>-18 4</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>17,-18,29.5,-18</points>
<connection>
<GID>99</GID>
<name>IN_2</name></connection>
<intersection>17 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>17,-34,29.5,-34</points>
<connection>
<GID>103</GID>
<name>IN_2</name></connection>
<intersection>17 3</intersection>
<intersection>25 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>25,-50.5,25,-34</points>
<intersection>-50.5 8</intersection>
<intersection>-34 6</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>25,-50.5,29.5,-50.5</points>
<connection>
<GID>107</GID>
<name>IN_2</name></connection>
<intersection>25 7</intersection></hsegment></shape></wire></page 3>
<page 4>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>54.5,-4</position>
<gparam>LABEL_TEXT DECODERS  (3*8)</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>BE_DECODER_3x8</type>
<position>46.5,-21.5</position>
<input>
<ID>ENABLE</ID>28 </input>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>30 </input>
<input>
<ID>IN_2</ID>29 </input>
<output>
<ID>OUT_0</ID>39 </output>
<output>
<ID>OUT_1</ID>38 </output>
<output>
<ID>OUT_2</ID>37 </output>
<output>
<ID>OUT_3</ID>36 </output>
<output>
<ID>OUT_4</ID>35 </output>
<output>
<ID>OUT_5</ID>34 </output>
<output>
<ID>OUT_6</ID>33 </output>
<output>
<ID>OUT_7</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_TOGGLE</type>
<position>17.5,-15.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_TOGGLE</type>
<position>17.5,-23.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>80</ID>
<type>AA_TOGGLE</type>
<position>17.5,-31.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>84</ID>
<type>AA_TOGGLE</type>
<position>17,-39.5</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>88</ID>
<type>GA_LED</type>
<position>63.5,-15.5</position>
<input>
<ID>N_in0</ID>32 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>GA_LED</type>
<position>63.5,-19.5</position>
<input>
<ID>N_in0</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>GA_LED</type>
<position>64,-24</position>
<input>
<ID>N_in0</ID>34 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>100</ID>
<type>GA_LED</type>
<position>64,-28</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>GA_LED</type>
<position>64,-32.5</position>
<input>
<ID>N_in0</ID>36 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>GA_LED</type>
<position>64.5,-36.5</position>
<input>
<ID>N_in0</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>GA_LED</type>
<position>64.5,-41</position>
<input>
<ID>N_in0</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>GA_LED</type>
<position>65,-45</position>
<input>
<ID>N_in0</ID>39 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-18,31.5,-15.5</points>
<intersection>-18 1</intersection>
<intersection>-15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-18,43.5,-18</points>
<connection>
<GID>73</GID>
<name>ENABLE</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-15.5,31.5,-15.5</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-23.5,31.5,-23</points>
<intersection>-23.5 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-23,43.5,-23</points>
<connection>
<GID>73</GID>
<name>IN_2</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-23.5,31.5,-23.5</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-31.5,31.5,-24</points>
<intersection>-31.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-24,43.5,-24</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-31.5,31.5,-31.5</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-39.5,34.5,-25</points>
<intersection>-39.5 2</intersection>
<intersection>-25 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-25,43.5,-25</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,-39.5,34.5,-39.5</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-18,56,-15.5</points>
<intersection>-18 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-15.5,62.5,-15.5</points>
<connection>
<GID>88</GID>
<name>N_in0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-18,56,-18</points>
<connection>
<GID>73</GID>
<name>OUT_7</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-19.5,56,-19</points>
<intersection>-19.5 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-19.5,62.5,-19.5</points>
<connection>
<GID>92</GID>
<name>N_in0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-19,56,-19</points>
<connection>
<GID>73</GID>
<name>OUT_6</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-24,56,-20</points>
<intersection>-24 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-24,63,-24</points>
<connection>
<GID>96</GID>
<name>N_in0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-20,56,-20</points>
<connection>
<GID>73</GID>
<name>OUT_5</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-28,55,-21</points>
<intersection>-28 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-28,63,-28</points>
<connection>
<GID>100</GID>
<name>N_in0</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-21,55,-21</points>
<connection>
<GID>73</GID>
<name>OUT_4</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-32.5,53.5,-22</points>
<intersection>-32.5 1</intersection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53.5,-32.5,63,-32.5</points>
<connection>
<GID>104</GID>
<name>N_in0</name></connection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-22,53.5,-22</points>
<connection>
<GID>73</GID>
<name>OUT_3</name></connection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-36.5,52.5,-23</points>
<intersection>-36.5 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-36.5,63.5,-36.5</points>
<connection>
<GID>108</GID>
<name>N_in0</name></connection>
<intersection>52.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-23,52.5,-23</points>
<connection>
<GID>73</GID>
<name>OUT_2</name></connection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51.5,-41,51.5,-24</points>
<intersection>-41 1</intersection>
<intersection>-24 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51.5,-41,63.5,-41</points>
<connection>
<GID>112</GID>
<name>N_in0</name></connection>
<intersection>51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-24,51.5,-24</points>
<connection>
<GID>73</GID>
<name>OUT_1</name></connection>
<intersection>51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-45,50.5,-25</points>
<intersection>-45 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-45,64,-45</points>
<connection>
<GID>116</GID>
<name>N_in0</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-25,50.5,-25</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire></page 4>
<page 5>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>62,-2.5</position>
<gparam>LABEL_TEXT ENCODERS    (8*3)</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_TOGGLE</type>
<position>14,-12</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_TOGGLE</type>
<position>14,-17.5</position>
<output>
<ID>OUT_0</ID>65 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_TOGGLE</type>
<position>14,-22</position>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_TOGGLE</type>
<position>14,-26.5</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>128</ID>
<type>AA_TOGGLE</type>
<position>14,-31.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_TOGGLE</type>
<position>14,-36</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_TOGGLE</type>
<position>14,-40.5</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_TOGGLE</type>
<position>14,-45</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>78.5,-16.5</position>
<input>
<ID>N_in0</ID>63 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>GA_LED</type>
<position>78.5,-30.5</position>
<input>
<ID>N_in0</ID>64 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>GA_LED</type>
<position>79,-46</position>
<input>
<ID>N_in0</ID>66 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>AE_OR4</type>
<position>51.5,-15</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>58 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>60 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>162</ID>
<type>AE_OR4</type>
<position>51.5,-28</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>62 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>60 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>164</ID>
<type>AE_OR4</type>
<position>52.5,-43.5</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>62 </input>
<input>
<ID>IN_2</ID>58 </input>
<input>
<ID>IN_3</ID>60 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>166</ID>
<type>AA_LABEL</type>
<position>96.5,-45.5</position>
<gparam>LABEL_TEXT Z=D1+D3+D5+D7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AA_LABEL</type>
<position>96,-16</position>
<gparam>LABEL_TEXT X=D4+D5+D6+D7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_LABEL</type>
<position>96.5,-30</position>
<gparam>LABEL_TEXT Y=D2+D3+D6+D7</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-31.5,20.5,-12</points>
<intersection>-31.5 2</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-12,48.5,-12</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-31.5,20.5,-31.5</points>
<connection>
<GID>128</GID>
<name>OUT_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-44.5,22.5,-14</points>
<intersection>-44.5 3</intersection>
<intersection>-36 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-14,48.5,-14</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-36,22.5,-36</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>22.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>22.5,-44.5,49.5,-44.5</points>
<connection>
<GID>164</GID>
<name>IN_2</name></connection>
<intersection>22.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-40.5,24,-16</points>
<intersection>-40.5 2</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24,-16,48.5,-16</points>
<connection>
<GID>160</GID>
<name>IN_2</name></connection>
<intersection>24 0</intersection>
<intersection>39 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-40.5,24,-40.5</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>24 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>39,-29,39,-16</points>
<intersection>-29 4</intersection>
<intersection>-16 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>39,-29,48.5,-29</points>
<connection>
<GID>162</GID>
<name>IN_2</name></connection>
<intersection>39 3</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-45,26,-18</points>
<intersection>-45 2</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-18,48.5,-18</points>
<connection>
<GID>160</GID>
<name>IN_3</name></connection>
<intersection>26 0</intersection>
<intersection>43 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-45,26,-45</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>26 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>43,-46.5,43,-18</points>
<intersection>-46.5 6</intersection>
<intersection>-31 4</intersection>
<intersection>-18 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>43,-31,48.5,-31</points>
<connection>
<GID>162</GID>
<name>IN_3</name></connection>
<intersection>43 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>43,-46.5,49.5,-46.5</points>
<connection>
<GID>164</GID>
<name>IN_3</name></connection>
<intersection>43 3</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-25,32,-22</points>
<intersection>-25 1</intersection>
<intersection>-22 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-25,48.5,-25</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-22,32,-22</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-27,32,-26.5</points>
<intersection>-27 1</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-27,48.5,-27</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<intersection>32 0</intersection>
<intersection>37 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>16,-26.5,32,-26.5</points>
<connection>
<GID>126</GID>
<name>OUT_0</name></connection>
<intersection>32 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37,-42.5,37,-27</points>
<intersection>-42.5 4</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37,-42.5,49.5,-42.5</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>37 3</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-16.5,66.5,-15</points>
<intersection>-16.5 1</intersection>
<intersection>-15 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-16.5,77.5,-16.5</points>
<connection>
<GID>154</GID>
<name>N_in0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-15,66.5,-15</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-30.5,66.5,-28</points>
<intersection>-30.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-30.5,77.5,-30.5</points>
<connection>
<GID>156</GID>
<name>N_in0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-28,66.5,-28</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32.5,-40.5,32.5,-10.5</points>
<intersection>-40.5 1</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32.5,-40.5,49.5,-40.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18,-10.5,32.5,-10.5</points>
<intersection>18 3</intersection>
<intersection>32.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>18,-17.5,18,-10.5</points>
<intersection>-17.5 4</intersection>
<intersection>-10.5 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>16,-17.5,18,-17.5</points>
<connection>
<GID>122</GID>
<name>OUT_0</name></connection>
<intersection>18 3</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-46,67,-43.5</points>
<intersection>-46 1</intersection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-46,78,-46</points>
<connection>
<GID>158</GID>
<name>N_in0</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-43.5,67,-43.5</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire></page 5>
<page 6>
<PageViewport>0,-3,122.4,-63.5</PageViewport>
<gate>
<ID>194</ID>
<type>AA_INVERTER</type>
<position>22,-17.5</position>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_INVERTER</type>
<position>22,-35.5</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>198</ID>
<type>AA_AND3</type>
<position>50,-56.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>68 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>59.5,-5.5</position>
<gparam>LABEL_TEXT DEMULTIPLEXERS   (1*4)</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_TOGGLE</type>
<position>12.5,-17.5</position>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_TOGGLE</type>
<position>13,-35.5</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>178</ID>
<type>GA_LED</type>
<position>83,-17.5</position>
<input>
<ID>N_in0</ID>77 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>GA_LED</type>
<position>83.5,-28.5</position>
<input>
<ID>N_in0</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>182</ID>
<type>GA_LED</type>
<position>83.5,-37.5</position>
<input>
<ID>N_in0</ID>75 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>GA_LED</type>
<position>84,-48.5</position>
<input>
<ID>N_in0</ID>74 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_TOGGLE</type>
<position>8,-48</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_AND3</type>
<position>48,-17</position>
<input>
<ID>IN_0</ID>69 </input>
<input>
<ID>IN_1</ID>70 </input>
<input>
<ID>IN_2</ID>68 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_AND3</type>
<position>48.5,-32.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>69 </input>
<input>
<ID>IN_2</ID>68 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_AND3</type>
<position>48,-46</position>
<input>
<ID>IN_0</ID>70 </input>
<input>
<ID>IN_1</ID>72 </input>
<input>
<ID>IN_2</ID>68 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29.5,-58.5,29.5,-19</points>
<intersection>-58.5 11</intersection>
<intersection>-48 1</intersection>
<intersection>-34.5 4</intersection>
<intersection>-19 6</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-48,45,-48</points>
<connection>
<GID>192</GID>
<name>IN_2</name></connection>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>29.5,-34.5,45.5,-34.5</points>
<connection>
<GID>190</GID>
<name>IN_2</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>29.5,-19,45,-19</points>
<connection>
<GID>188</GID>
<name>IN_2</name></connection>
<intersection>29.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>29.5,-58.5,47,-58.5</points>
<connection>
<GID>198</GID>
<name>IN_2</name></connection>
<intersection>29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-27,45,-27</points>
<intersection>15 5</intersection>
<intersection>19 4</intersection>
<intersection>40.5 3</intersection>
<intersection>45 7</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>40.5,-32.5,40.5,-27</points>
<intersection>-32.5 6</intersection>
<intersection>-27 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>19,-35.5,19,-27</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>-27 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>15,-35.5,15,-27</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>40.5,-32.5,45.5,-32.5</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>40.5 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>45,-27,45,-15</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>-27 1</intersection></vsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>14.5,-12,37.5,-12</points>
<intersection>14.5 6</intersection>
<intersection>19 5</intersection>
<intersection>37.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37.5,-44,37.5,-12</points>
<intersection>-44 4</intersection>
<intersection>-17 7</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37.5,-44,45,-44</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>37.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>19,-17.5,19,-12</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>-12 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>14.5,-17.5,14.5,-12</points>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>37.5,-17,45,-17</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<intersection>37.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-56.5,25.5,-35.5</points>
<intersection>-56.5 1</intersection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-56.5,47,-56.5</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>25.5 0</intersection>
<intersection>40 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-35.5,25.5,-35.5</points>
<connection>
<GID>196</GID>
<name>OUT_0</name></connection>
<intersection>25.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>40,-56.5,40,-46</points>
<intersection>-56.5 1</intersection>
<intersection>-46 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>40,-46,45,-46</points>
<connection>
<GID>192</GID>
<name>IN_1</name></connection>
<intersection>40 3</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28,-54.5,28,-17.5</points>
<intersection>-54.5 2</intersection>
<intersection>-30.5 3</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-17.5,28,-17.5</points>
<connection>
<GID>194</GID>
<name>OUT_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-54.5,47,-54.5</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>28,-30.5,45.5,-30.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>28 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-56.5,68,-48.5</points>
<intersection>-56.5 2</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-48.5,83,-48.5</points>
<connection>
<GID>184</GID>
<name>N_in0</name></connection>
<intersection>68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>53,-56.5,68,-56.5</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-46,66.5,-37.5</points>
<intersection>-46 2</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-37.5,82.5,-37.5</points>
<connection>
<GID>182</GID>
<name>N_in0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-46,66.5,-46</points>
<connection>
<GID>192</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-32.5,67,-28.5</points>
<intersection>-32.5 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67,-28.5,82.5,-28.5</points>
<connection>
<GID>180</GID>
<name>N_in0</name></connection>
<intersection>67 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51.5,-32.5,67,-32.5</points>
<connection>
<GID>190</GID>
<name>OUT</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-17.5,66.5,-17</points>
<intersection>-17.5 1</intersection>
<intersection>-17 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-17.5,82,-17.5</points>
<connection>
<GID>178</GID>
<name>N_in0</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-17,66.5,-17</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire></page 6>
<page 7>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport>
<gate>
<ID>200</ID>
<type>AA_LABEL</type>
<position>60,-3.5</position>
<gparam>LABEL_TEXT MULTIPLEXERS   (4*1)</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>AA_TOGGLE</type>
<position>18,-13.5</position>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>204</ID>
<type>AA_TOGGLE</type>
<position>18.5,-21.5</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>206</ID>
<type>AA_TOGGLE</type>
<position>18,-29</position>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>208</ID>
<type>AA_TOGGLE</type>
<position>18,-37</position>
<output>
<ID>OUT_0</ID>81 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>210</ID>
<type>GA_LED</type>
<position>95.5,-24.5</position>
<input>
<ID>N_in0</ID>93 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>212</ID>
<type>AA_AND3</type>
<position>52,-13.5</position>
<input>
<ID>IN_0</ID>78 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>83 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_AND3</type>
<position>52,-25</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>83 </input>
<input>
<ID>IN_2</ID>84 </input>
<output>
<ID>OUT</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_AND3</type>
<position>52.5,-35.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>85 </input>
<input>
<ID>IN_2</ID>82 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_AND3</type>
<position>52.5,-44.5</position>
<input>
<ID>IN_0</ID>81 </input>
<input>
<ID>IN_1</ID>84 </input>
<input>
<ID>IN_2</ID>85 </input>
<output>
<ID>OUT</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_TOGGLE</type>
<position>18.5,-44.5</position>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_TOGGLE</type>
<position>18.5,-50</position>
<output>
<ID>OUT_0</ID>83 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>224</ID>
<type>AA_INVERTER</type>
<position>27.5,-43.5</position>
<input>
<ID>IN_0</ID>82 </input>
<output>
<ID>OUT_0</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>226</ID>
<type>AA_INVERTER</type>
<position>28,-50</position>
<input>
<ID>IN_0</ID>83 </input>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>228</ID>
<type>AE_OR4</type>
<position>75,-23</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>90 </input>
<input>
<ID>IN_2</ID>91 </input>
<input>
<ID>IN_3</ID>92 </input>
<output>
<ID>OUT</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-13.5,34.5,-11.5</points>
<intersection>-13.5 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-11.5,49,-11.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,-13.5,34.5,-13.5</points>
<connection>
<GID>202</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-23,34.5,-21.5</points>
<intersection>-23 1</intersection>
<intersection>-21.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-23,49,-23</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20.5,-21.5,34.5,-21.5</points>
<connection>
<GID>204</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-33.5,34.5,-29</points>
<intersection>-33.5 1</intersection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-33.5,49.5,-33.5</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,-29,34.5,-29</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34.5,-42.5,34.5,-37</points>
<intersection>-42.5 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34.5,-42.5,49.5,-42.5</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>34.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20,-37,34.5,-37</points>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection>
<intersection>34.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-44.5,22.5,-40</points>
<intersection>-44.5 2</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-40,46,-40</points>
<intersection>22.5 0</intersection>
<intersection>24.5 5</intersection>
<intersection>46 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20.5,-44.5,22.5,-44.5</points>
<connection>
<GID>220</GID>
<name>OUT_0</name></connection>
<intersection>22.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>46,-40,46,-37.5</points>
<intersection>-40 1</intersection>
<intersection>-37.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36.5,-37.5,49.5,-37.5</points>
<connection>
<GID>216</GID>
<name>IN_2</name></connection>
<intersection>36.5 6</intersection>
<intersection>46 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>24.5,-43.5,24.5,-40</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>-40 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>36.5,-37.5,36.5,-13.5</points>
<intersection>-37.5 4</intersection>
<intersection>-13.5 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>36.5,-13.5,49,-13.5</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<intersection>36.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-54,45,-54</points>
<intersection>20.5 8</intersection>
<intersection>25 7</intersection>
<intersection>45 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>45,-54,45,-15.5</points>
<intersection>-54 1</intersection>
<intersection>-25 4</intersection>
<intersection>-15.5 6</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>45,-25,49,-25</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>45 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>45,-15.5,49,-15.5</points>
<connection>
<GID>212</GID>
<name>IN_2</name></connection>
<intersection>45 3</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>25,-54,25,-50</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>-54 1</intersection></vsegment>
<vsegment>
<ID>8</ID>
<points>20.5,-54,20.5,-50</points>
<connection>
<GID>222</GID>
<name>OUT_0</name></connection>
<intersection>-54 1</intersection></vsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-44.5,40,-43.5</points>
<intersection>-44.5 1</intersection>
<intersection>-43.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-44.5,49.5,-44.5</points>
<connection>
<GID>218</GID>
<name>IN_1</name></connection>
<intersection>40 0</intersection>
<intersection>47.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-43.5,40,-43.5</points>
<connection>
<GID>224</GID>
<name>OUT_0</name></connection>
<intersection>40 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47.5,-44.5,47.5,-27</points>
<intersection>-44.5 1</intersection>
<intersection>-27 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>47.5,-27,49,-27</points>
<connection>
<GID>214</GID>
<name>IN_2</name></connection>
<intersection>47.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-50,40,-46.5</points>
<intersection>-50 2</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40,-46.5,49.5,-46.5</points>
<connection>
<GID>218</GID>
<name>IN_2</name></connection>
<intersection>40 0</intersection>
<intersection>42.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-50,40,-50</points>
<connection>
<GID>226</GID>
<name>OUT_0</name></connection>
<intersection>40 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>42.5,-46.5,42.5,-35.5</points>
<intersection>-46.5 1</intersection>
<intersection>-35.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>42.5,-35.5,49.5,-35.5</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<intersection>42.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-20,63.5,-13.5</points>
<intersection>-20 1</intersection>
<intersection>-13.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-20,72,-20</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55,-13.5,63.5,-13.5</points>
<connection>
<GID>212</GID>
<name>OUT</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-25,63.5,-22</points>
<intersection>-25 2</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-22,72,-22</points>
<connection>
<GID>228</GID>
<name>IN_1</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55,-25,63.5,-25</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>64.5,-35.5,64.5,-24</points>
<intersection>-35.5 2</intersection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64.5,-24,72,-24</points>
<connection>
<GID>228</GID>
<name>IN_2</name></connection>
<intersection>64.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-35.5,64.5,-35.5</points>
<connection>
<GID>216</GID>
<name>OUT</name></connection>
<intersection>64.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-44.5,66.5,-26</points>
<intersection>-44.5 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66.5,-26,72,-26</points>
<connection>
<GID>228</GID>
<name>IN_3</name></connection>
<intersection>66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-44.5,66.5,-44.5</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<intersection>66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-24.5,86.5,-23</points>
<intersection>-24.5 1</intersection>
<intersection>-23 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-24.5,94.5,-24.5</points>
<connection>
<GID>210</GID>
<name>N_in0</name></connection>
<intersection>86.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>79,-23,86.5,-23</points>
<connection>
<GID>228</GID>
<name>OUT</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire></page 7>
<page 8>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>58,-3.5</position>
<gparam>LABEL_TEXT MULTIPLEXERS  (4*1)</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AE_MUX_4x1</type>
<position>52.5,-28</position>
<input>
<ID>IN_0</ID>67 </input>
<input>
<ID>IN_1</ID>54 </input>
<input>
<ID>IN_2</ID>41 </input>
<input>
<ID>IN_3</ID>40 </input>
<output>
<ID>OUT</ID>87 </output>
<input>
<ID>SEL_0</ID>86 </input>
<input>
<ID>SEL_1</ID>71 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_TOGGLE</type>
<position>15,-19</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_TOGGLE</type>
<position>15,-26</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_TOGGLE</type>
<position>15,-33.5</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_TOGGLE</type>
<position>15,-40.5</position>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>78</ID>
<type>AA_TOGGLE</type>
<position>47.5,-13.5</position>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_TOGGLE</type>
<position>53,-12.5</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>94</ID>
<type>GA_LED</type>
<position>68,-27</position>
<input>
<ID>N_in0</ID>87 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-25,33,-19</points>
<intersection>-25 1</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-25,49.5,-25</points>
<connection>
<GID>53</GID>
<name>IN_3</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-19,33,-19</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-27,33,-26</points>
<intersection>-27 1</intersection>
<intersection>-26 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-27,49.5,-27</points>
<connection>
<GID>53</GID>
<name>IN_2</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-26,33,-26</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-33.5,33,-29</points>
<intersection>-33.5 2</intersection>
<intersection>-29 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-29,49.5,-29</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-33.5,33,-33.5</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-40.5,35.5,-31</points>
<intersection>-40.5 2</intersection>
<intersection>-31 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35.5,-31,49.5,-31</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>35.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>17,-40.5,35.5,-40.5</points>
<connection>
<GID>74</GID>
<name>OUT_0</name></connection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>52.5,-23,52.5,-18.5</points>
<connection>
<GID>53</GID>
<name>SEL_1</name></connection>
<intersection>-18.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>47.5,-18.5,47.5,-15.5</points>
<connection>
<GID>78</GID>
<name>OUT_0</name></connection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>47.5,-18.5,52.5,-18.5</points>
<intersection>47.5 1</intersection>
<intersection>52.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-23,53.5,-18.5</points>
<connection>
<GID>53</GID>
<name>SEL_0</name></connection>
<intersection>-18.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>53,-18.5,53,-14.5</points>
<connection>
<GID>86</GID>
<name>OUT_0</name></connection>
<intersection>-18.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>53,-18.5,53.5,-18.5</points>
<intersection>53 1</intersection>
<intersection>53.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-28,61,-27</points>
<intersection>-28 2</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-27,67,-27</points>
<connection>
<GID>94</GID>
<name>N_in0</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55.5,-28,61,-28</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire></page 8>
<page 9>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>53,-3.5</position>
<gparam>LABEL_TEXT D FLIP FLOP</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>BA_NAND2</type>
<position>32.5,-18</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>BA_NAND2</type>
<position>45.5,-37.5</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>121</ID>
<type>BA_NAND2</type>
<position>30,-38</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>125</ID>
<type>BB_CLOCK</type>
<position>7.5,-24.5</position>
<output>
<ID>CLK</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_TOGGLE</type>
<position>7.5,-12.5</position>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>136</ID>
<type>BA_NAND2</type>
<position>63,-38.5</position>
<input>
<ID>IN_0</ID>101 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>BA_NAND2</type>
<position>57,-16</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>99 </input>
<output>
<ID>OUT</ID>100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>140</ID>
<type>GA_LED</type>
<position>76,-16.5</position>
<input>
<ID>N_in0</ID>100 </input>
<input>
<ID>N_in1</ID>101 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>142</ID>
<type>GA_LED</type>
<position>81,-38</position>
<input>
<ID>N_in0</ID>99 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>AA_LABEL</type>
<position>83,-15.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>146</ID>
<type>AA_LABEL</type>
<position>87.5,-37.5</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-30.5,20.5,-19</points>
<intersection>-30.5 3</intersection>
<intersection>-24.5 2</intersection>
<intersection>-19 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-19,29.5,-19</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11.5,-24.5,20.5,-24.5</points>
<connection>
<GID>125</GID>
<name>CLK</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>20.5,-30.5,42.5,-30.5</points>
<intersection>20.5 0</intersection>
<intersection>27 5</intersection>
<intersection>42.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>42.5,-36.5,42.5,-30.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>-30.5 3</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>27,-37,27,-30.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>-30.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-17,19.5,-12.5</points>
<intersection>-17 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-17,29.5,-17</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>13.5 3</intersection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>9.5,-12.5,19.5,-12.5</points>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<intersection>19.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13.5,-39,13.5,-17</points>
<intersection>-39 4</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>13.5,-39,27,-39</points>
<connection>
<GID>121</GID>
<name>IN_1</name></connection>
<intersection>13.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-38.5,37.5,-38</points>
<intersection>-38.5 1</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>37.5,-38.5,42.5,-38.5</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-38,37.5,-38</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-38,73,-27.5</points>
<intersection>-38 1</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-38,80,-38</points>
<connection>
<GID>142</GID>
<name>N_in0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54,-27.5,73,-27.5</points>
<intersection>54 3</intersection>
<intersection>67.5 4</intersection>
<intersection>73 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54,-27.5,54,-17</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>-27.5 2</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>67.5,-38.5,67.5,-27.5</points>
<intersection>-38.5 5</intersection>
<intersection>-27.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>66,-38.5,67.5,-38.5</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<intersection>67.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-16.5,67.5,-16</points>
<intersection>-16.5 1</intersection>
<intersection>-16 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>67.5,-16.5,75,-16.5</points>
<connection>
<GID>140</GID>
<name>N_in0</name></connection>
<intersection>67.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60,-16,67.5,-16</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-21.5,68.5,-16.5</points>
<intersection>-21.5 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68.5,-16.5,77,-16.5</points>
<connection>
<GID>140</GID>
<name>N_in1</name></connection>
<intersection>68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60,-21.5,68.5,-21.5</points>
<intersection>60 3</intersection>
<intersection>68.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>60,-37.5,60,-21.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-21.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>102</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-18,44.5,-15</points>
<intersection>-18 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-15,54,-15</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>35.5,-18,44.5,-18</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-39.5,54,-37.5</points>
<intersection>-39.5 1</intersection>
<intersection>-37.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-39.5,60,-39.5</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48.5,-37.5,54,-37.5</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire></page 9></circuit>